module player(input wire clk, input wire [5:0] i, input wire [7:0] j, output reg [2:0] pixel);
  (* rom_style = "block" *)

//signal declarations
  reg [5:0] row_reg;
  reg [7:0] col_reg;
  always @(posedge clk)
	begin
	row_reg <= i;
	col_reg <= j;
	end


always @*
    case ({row_reg, col_reg})
      14'b00000000000000: pixel[2:0] = 3'b000;
      14'b00000000000001: pixel[2:0] = 3'b000;
      14'b00000000000010: pixel[2:0] = 3'b000;
      14'b00000000000011: pixel[2:0] = 3'b000;
      14'b00000000000100: pixel[2:0] = 3'b000;
      14'b00000000000101: pixel[2:0] = 3'b000;
      14'b00000000000110: pixel[2:0] = 3'b000;
      14'b00000000000111: pixel[2:0] = 3'b000;
      14'b00000000001000: pixel[2:0] = 3'b000;
      14'b00000000001001: pixel[2:0] = 3'b000;
      14'b00000000001010: pixel[2:0] = 3'b000;
      14'b00000000001011: pixel[2:0] = 3'b000;
      14'b00000000001100: pixel[2:0] = 3'b000;
      14'b00000000001101: pixel[2:0] = 3'b000;
      14'b00000000001110: pixel[2:0] = 3'b000;
      14'b00000000001111: pixel[2:0] = 3'b000;
      14'b00000000010000: pixel[2:0] = 3'b000;
      14'b00000000010001: pixel[2:0] = 3'b000;
      14'b00000000010010: pixel[2:0] = 3'b000;
      14'b00000000010011: pixel[2:0] = 3'b000;
      14'b00000000010100: pixel[2:0] = 3'b000;
      14'b00000000010101: pixel[2:0] = 3'b000;
      14'b00000000010110: pixel[2:0] = 3'b000;
      14'b00000000010111: pixel[2:0] = 3'b000;
      14'b00000000011000: pixel[2:0] = 3'b000;
      14'b00000000011001: pixel[2:0] = 3'b000;
      14'b00000000011010: pixel[2:0] = 3'b000;
      14'b00000000011011: pixel[2:0] = 3'b000;
      14'b00000000011100: pixel[2:0] = 3'b000;
      14'b00000000011101: pixel[2:0] = 3'b000;
      14'b00000000011110: pixel[2:0] = 3'b000;
      14'b00000000011111: pixel[2:0] = 3'b000;
      14'b00000000100000: pixel[2:0] = 3'b000;
      14'b00000000100001: pixel[2:0] = 3'b000;
      14'b00000000100010: pixel[2:0] = 3'b000;
      14'b00000000100011: pixel[2:0] = 3'b000;
      14'b00000000100100: pixel[2:0] = 3'b000;
      14'b00000000100101: pixel[2:0] = 3'b000;
      14'b00000000100110: pixel[2:0] = 3'b000;
      14'b00000000100111: pixel[2:0] = 3'b000;
      14'b00000000101000: pixel[2:0] = 3'b000;
      14'b00000000101001: pixel[2:0] = 3'b000;
      14'b00000000101010: pixel[2:0] = 3'b000;
      14'b00000000101011: pixel[2:0] = 3'b000;
      14'b00000000101100: pixel[2:0] = 3'b000;
      14'b00000000101101: pixel[2:0] = 3'b000;
      14'b00000000101110: pixel[2:0] = 3'b000;
      14'b00000000101111: pixel[2:0] = 3'b000;
      14'b00000000110000: pixel[2:0] = 3'b000;
      14'b00000000110001: pixel[2:0] = 3'b000;
      14'b00000000110010: pixel[2:0] = 3'b000;
      14'b00000000110011: pixel[2:0] = 3'b000;
      14'b00000000110100: pixel[2:0] = 3'b000;
      14'b00000000110101: pixel[2:0] = 3'b000;
      14'b00000000110110: pixel[2:0] = 3'b000;
      14'b00000000110111: pixel[2:0] = 3'b000;
      14'b00000000111000: pixel[2:0] = 3'b000;
      14'b00000000111001: pixel[2:0] = 3'b000;
      14'b00000000111010: pixel[2:0] = 3'b000;
      14'b00000000111011: pixel[2:0] = 3'b000;
      14'b00000000111100: pixel[2:0] = 3'b000;
      14'b00000000111101: pixel[2:0] = 3'b000;
      14'b00000000111110: pixel[2:0] = 3'b000;
      14'b00000000111111: pixel[2:0] = 3'b000;
      14'b00000001000000: pixel[2:0] = 3'b000;
      14'b00000001000001: pixel[2:0] = 3'b000;
      14'b00000001000010: pixel[2:0] = 3'b000;
      14'b00000001000011: pixel[2:0] = 3'b000;
      14'b00000001000100: pixel[2:0] = 3'b000;
      14'b00000001000101: pixel[2:0] = 3'b000;
      14'b00000001000110: pixel[2:0] = 3'b000;
      14'b00000001000111: pixel[2:0] = 3'b000;
      14'b00000001001000: pixel[2:0] = 3'b000;
      14'b00000001001001: pixel[2:0] = 3'b000;
      14'b00000001001010: pixel[2:0] = 3'b000;
      14'b00000001001011: pixel[2:0] = 3'b000;
      14'b00000001001100: pixel[2:0] = 3'b000;
      14'b00000001001101: pixel[2:0] = 3'b000;
      14'b00000001001110: pixel[2:0] = 3'b000;
      14'b00000001001111: pixel[2:0] = 3'b000;
      14'b00000001010000: pixel[2:0] = 3'b000;
      14'b00000001010001: pixel[2:0] = 3'b000;
      14'b00000001010010: pixel[2:0] = 3'b000;
      14'b00000001010011: pixel[2:0] = 3'b000;
      14'b00000001010100: pixel[2:0] = 3'b000;
      14'b00000001010101: pixel[2:0] = 3'b000;
      14'b00000001010110: pixel[2:0] = 3'b000;
      14'b00000001010111: pixel[2:0] = 3'b000;
      14'b00000001011000: pixel[2:0] = 3'b000;
      14'b00000001011001: pixel[2:0] = 3'b000;
      14'b00000001011010: pixel[2:0] = 3'b000;
      14'b00000001011011: pixel[2:0] = 3'b000;
      14'b00000001011100: pixel[2:0] = 3'b000;
      14'b00000001011101: pixel[2:0] = 3'b000;
      14'b00000001011110: pixel[2:0] = 3'b000;
      14'b00000001011111: pixel[2:0] = 3'b000;
      14'b00000001100000: pixel[2:0] = 3'b000;
      14'b00000001100001: pixel[2:0] = 3'b000;
      14'b00000001100010: pixel[2:0] = 3'b000;
      14'b00000001100011: pixel[2:0] = 3'b000;
      14'b00000001100100: pixel[2:0] = 3'b000;
      14'b00000001100101: pixel[2:0] = 3'b000;
      14'b00000001100110: pixel[2:0] = 3'b000;
      14'b00000001100111: pixel[2:0] = 3'b000;
      14'b00000001101000: pixel[2:0] = 3'b000;
      14'b00000001101001: pixel[2:0] = 3'b000;
      14'b00000001101010: pixel[2:0] = 3'b000;
      14'b00000001101011: pixel[2:0] = 3'b000;
      14'b00000001101100: pixel[2:0] = 3'b000;
      14'b00000001101101: pixel[2:0] = 3'b000;
      14'b00000001101110: pixel[2:0] = 3'b000;
      14'b00000001101111: pixel[2:0] = 3'b000;
      14'b00000001110000: pixel[2:0] = 3'b000;
      14'b00000001110001: pixel[2:0] = 3'b000;
      14'b00000001110010: pixel[2:0] = 3'b000;
      14'b00000001110011: pixel[2:0] = 3'b000;
      14'b00000001110100: pixel[2:0] = 3'b000;
      14'b00000001110101: pixel[2:0] = 3'b000;
      14'b00000001110110: pixel[2:0] = 3'b000;
      14'b00000001110111: pixel[2:0] = 3'b000;
      14'b00000001111000: pixel[2:0] = 3'b000;
      14'b00000001111001: pixel[2:0] = 3'b000;
      14'b00000001111010: pixel[2:0] = 3'b000;
      14'b00000001111011: pixel[2:0] = 3'b000;
      14'b00000001111100: pixel[2:0] = 3'b000;
      14'b00000001111101: pixel[2:0] = 3'b000;
      14'b00000001111110: pixel[2:0] = 3'b000;
      14'b00000001111111: pixel[2:0] = 3'b000;
      14'b00000010000000: pixel[2:0] = 3'b000;
      14'b00000010000001: pixel[2:0] = 3'b000;
      14'b00000010000010: pixel[2:0] = 3'b000;
      14'b00000010000011: pixel[2:0] = 3'b000;
      14'b00000010000100: pixel[2:0] = 3'b000;
      14'b00000010000101: pixel[2:0] = 3'b000;
      14'b00000010000110: pixel[2:0] = 3'b000;
      14'b00000010000111: pixel[2:0] = 3'b000;
      14'b00000100000000: pixel[2:0] = 3'b000;
      14'b00000100000001: pixel[2:0] = 3'b000;
      14'b00000100000010: pixel[2:0] = 3'b000;
      14'b00000100000011: pixel[2:0] = 3'b000;
      14'b00000100000100: pixel[2:0] = 3'b000;
      14'b00000100000101: pixel[2:0] = 3'b000;
      14'b00000100000110: pixel[2:0] = 3'b000;
      14'b00000100000111: pixel[2:0] = 3'b000;
      14'b00000100001000: pixel[2:0] = 3'b000;
      14'b00000100001001: pixel[2:0] = 3'b000;
      14'b00000100001010: pixel[2:0] = 3'b000;
      14'b00000100001011: pixel[2:0] = 3'b000;
      14'b00000100001100: pixel[2:0] = 3'b000;
      14'b00000100001101: pixel[2:0] = 3'b000;
      14'b00000100001110: pixel[2:0] = 3'b000;
      14'b00000100001111: pixel[2:0] = 3'b000;
      14'b00000100010000: pixel[2:0] = 3'b000;
      14'b00000100010001: pixel[2:0] = 3'b000;
      14'b00000100010010: pixel[2:0] = 3'b000;
      14'b00000100010011: pixel[2:0] = 3'b000;
      14'b00000100010100: pixel[2:0] = 3'b000;
      14'b00000100010101: pixel[2:0] = 3'b000;
      14'b00000100010110: pixel[2:0] = 3'b000;
      14'b00000100010111: pixel[2:0] = 3'b000;
      14'b00000100011000: pixel[2:0] = 3'b000;
      14'b00000100011001: pixel[2:0] = 3'b000;
      14'b00000100011010: pixel[2:0] = 3'b000;
      14'b00000100011011: pixel[2:0] = 3'b000;
      14'b00000100011100: pixel[2:0] = 3'b000;
      14'b00000100011101: pixel[2:0] = 3'b000;
      14'b00000100011110: pixel[2:0] = 3'b000;
      14'b00000100011111: pixel[2:0] = 3'b000;
      14'b00000100100000: pixel[2:0] = 3'b000;
      14'b00000100100001: pixel[2:0] = 3'b000;
      14'b00000100100010: pixel[2:0] = 3'b000;
      14'b00000100100011: pixel[2:0] = 3'b000;
      14'b00000100100100: pixel[2:0] = 3'b000;
      14'b00000100100101: pixel[2:0] = 3'b000;
      14'b00000100100110: pixel[2:0] = 3'b000;
      14'b00000100100111: pixel[2:0] = 3'b000;
      14'b00000100101000: pixel[2:0] = 3'b000;
      14'b00000100101001: pixel[2:0] = 3'b000;
      14'b00000100101010: pixel[2:0] = 3'b000;
      14'b00000100101011: pixel[2:0] = 3'b000;
      14'b00000100101100: pixel[2:0] = 3'b000;
      14'b00000100101101: pixel[2:0] = 3'b000;
      14'b00000100101110: pixel[2:0] = 3'b000;
      14'b00000100101111: pixel[2:0] = 3'b000;
      14'b00000100110000: pixel[2:0] = 3'b000;
      14'b00000100110001: pixel[2:0] = 3'b000;
      14'b00000100110010: pixel[2:0] = 3'b000;
      14'b00000100110011: pixel[2:0] = 3'b000;
      14'b00000100110100: pixel[2:0] = 3'b000;
      14'b00000100110101: pixel[2:0] = 3'b000;
      14'b00000100110110: pixel[2:0] = 3'b000;
      14'b00000100110111: pixel[2:0] = 3'b000;
      14'b00000100111000: pixel[2:0] = 3'b000;
      14'b00000100111001: pixel[2:0] = 3'b000;
      14'b00000100111010: pixel[2:0] = 3'b000;
      14'b00000100111011: pixel[2:0] = 3'b000;
      14'b00000100111100: pixel[2:0] = 3'b000;
      14'b00000100111101: pixel[2:0] = 3'b000;
      14'b00000100111110: pixel[2:0] = 3'b000;
      14'b00000100111111: pixel[2:0] = 3'b000;
      14'b00000101000000: pixel[2:0] = 3'b000;
      14'b00000101000001: pixel[2:0] = 3'b000;
      14'b00000101000010: pixel[2:0] = 3'b000;
      14'b00000101000011: pixel[2:0] = 3'b000;
      14'b00000101000100: pixel[2:0] = 3'b000;
      14'b00000101000101: pixel[2:0] = 3'b000;
      14'b00000101000110: pixel[2:0] = 3'b000;
      14'b00000101000111: pixel[2:0] = 3'b000;
      14'b00000101001000: pixel[2:0] = 3'b000;
      14'b00000101001001: pixel[2:0] = 3'b000;
      14'b00000101001010: pixel[2:0] = 3'b000;
      14'b00000101001011: pixel[2:0] = 3'b000;
      14'b00000101001100: pixel[2:0] = 3'b000;
      14'b00000101001101: pixel[2:0] = 3'b000;
      14'b00000101001110: pixel[2:0] = 3'b000;
      14'b00000101001111: pixel[2:0] = 3'b000;
      14'b00000101010000: pixel[2:0] = 3'b000;
      14'b00000101010001: pixel[2:0] = 3'b000;
      14'b00000101010010: pixel[2:0] = 3'b000;
      14'b00000101010011: pixel[2:0] = 3'b000;
      14'b00000101010100: pixel[2:0] = 3'b000;
      14'b00000101010101: pixel[2:0] = 3'b000;
      14'b00000101010110: pixel[2:0] = 3'b000;
      14'b00000101010111: pixel[2:0] = 3'b000;
      14'b00000101011000: pixel[2:0] = 3'b000;
      14'b00000101011001: pixel[2:0] = 3'b000;
      14'b00000101011010: pixel[2:0] = 3'b000;
      14'b00000101011011: pixel[2:0] = 3'b000;
      14'b00000101011100: pixel[2:0] = 3'b000;
      14'b00000101011101: pixel[2:0] = 3'b000;
      14'b00000101011110: pixel[2:0] = 3'b000;
      14'b00000101011111: pixel[2:0] = 3'b000;
      14'b00000101100000: pixel[2:0] = 3'b000;
      14'b00000101100001: pixel[2:0] = 3'b000;
      14'b00000101100010: pixel[2:0] = 3'b000;
      14'b00000101100011: pixel[2:0] = 3'b000;
      14'b00000101100100: pixel[2:0] = 3'b000;
      14'b00000101100101: pixel[2:0] = 3'b000;
      14'b00000101100110: pixel[2:0] = 3'b000;
      14'b00000101100111: pixel[2:0] = 3'b000;
      14'b00000101101000: pixel[2:0] = 3'b000;
      14'b00000101101001: pixel[2:0] = 3'b000;
      14'b00000101101010: pixel[2:0] = 3'b000;
      14'b00000101101011: pixel[2:0] = 3'b000;
      14'b00000101101100: pixel[2:0] = 3'b000;
      14'b00000101101101: pixel[2:0] = 3'b000;
      14'b00000101101110: pixel[2:0] = 3'b000;
      14'b00000101101111: pixel[2:0] = 3'b000;
      14'b00000101110000: pixel[2:0] = 3'b000;
      14'b00000101110001: pixel[2:0] = 3'b000;
      14'b00000101110010: pixel[2:0] = 3'b000;
      14'b00000101110011: pixel[2:0] = 3'b000;
      14'b00000101110100: pixel[2:0] = 3'b000;
      14'b00000101110101: pixel[2:0] = 3'b000;
      14'b00000101110110: pixel[2:0] = 3'b000;
      14'b00000101110111: pixel[2:0] = 3'b000;
      14'b00000101111000: pixel[2:0] = 3'b000;
      14'b00000101111001: pixel[2:0] = 3'b000;
      14'b00000101111010: pixel[2:0] = 3'b000;
      14'b00000101111011: pixel[2:0] = 3'b000;
      14'b00000101111100: pixel[2:0] = 3'b000;
      14'b00000101111101: pixel[2:0] = 3'b000;
      14'b00000101111110: pixel[2:0] = 3'b000;
      14'b00000101111111: pixel[2:0] = 3'b000;
      14'b00000110000000: pixel[2:0] = 3'b000;
      14'b00000110000001: pixel[2:0] = 3'b000;
      14'b00000110000010: pixel[2:0] = 3'b000;
      14'b00000110000011: pixel[2:0] = 3'b000;
      14'b00000110000100: pixel[2:0] = 3'b000;
      14'b00000110000101: pixel[2:0] = 3'b000;
      14'b00000110000110: pixel[2:0] = 3'b000;
      14'b00000110000111: pixel[2:0] = 3'b000;
      14'b00001000000000: pixel[2:0] = 3'b000;
      14'b00001000000001: pixel[2:0] = 3'b000;
      14'b00001000000010: pixel[2:0] = 3'b111;
      14'b00001000000011: pixel[2:0] = 3'b111;
      14'b00001000000100: pixel[2:0] = 3'b111;
      14'b00001000000101: pixel[2:0] = 3'b111;
      14'b00001000000110: pixel[2:0] = 3'b111;
      14'b00001000000111: pixel[2:0] = 3'b111;
      14'b00001000001000: pixel[2:0] = 3'b111;
      14'b00001000001001: pixel[2:0] = 3'b111;
      14'b00001000001010: pixel[2:0] = 3'b111;
      14'b00001000001011: pixel[2:0] = 3'b111;
      14'b00001000001100: pixel[2:0] = 3'b111;
      14'b00001000001101: pixel[2:0] = 3'b000;
      14'b00001000001110: pixel[2:0] = 3'b000;
      14'b00001000001111: pixel[2:0] = 3'b000;
      14'b00001000010000: pixel[2:0] = 3'b000;
      14'b00001000010001: pixel[2:0] = 3'b000;
      14'b00001000010010: pixel[2:0] = 3'b000;
      14'b00001000010011: pixel[2:0] = 3'b000;
      14'b00001000010100: pixel[2:0] = 3'b000;
      14'b00001000010101: pixel[2:0] = 3'b000;
      14'b00001000010110: pixel[2:0] = 3'b000;
      14'b00001000010111: pixel[2:0] = 3'b000;
      14'b00001000011000: pixel[2:0] = 3'b000;
      14'b00001000011001: pixel[2:0] = 3'b111;
      14'b00001000011010: pixel[2:0] = 3'b111;
      14'b00001000011011: pixel[2:0] = 3'b111;
      14'b00001000011100: pixel[2:0] = 3'b111;
      14'b00001000011101: pixel[2:0] = 3'b111;
      14'b00001000011110: pixel[2:0] = 3'b000;
      14'b00001000011111: pixel[2:0] = 3'b000;
      14'b00001000100000: pixel[2:0] = 3'b000;
      14'b00001000100001: pixel[2:0] = 3'b000;
      14'b00001000100010: pixel[2:0] = 3'b000;
      14'b00001000100011: pixel[2:0] = 3'b000;
      14'b00001000100100: pixel[2:0] = 3'b000;
      14'b00001000100101: pixel[2:0] = 3'b000;
      14'b00001000100110: pixel[2:0] = 3'b000;
      14'b00001000100111: pixel[2:0] = 3'b000;
      14'b00001000101000: pixel[2:0] = 3'b000;
      14'b00001000101001: pixel[2:0] = 3'b000;
      14'b00001000101010: pixel[2:0] = 3'b000;
      14'b00001000101011: pixel[2:0] = 3'b000;
      14'b00001000101100: pixel[2:0] = 3'b000;
      14'b00001000101101: pixel[2:0] = 3'b000;
      14'b00001000101110: pixel[2:0] = 3'b000;
      14'b00001000101111: pixel[2:0] = 3'b000;
      14'b00001000110000: pixel[2:0] = 3'b000;
      14'b00001000110001: pixel[2:0] = 3'b000;
      14'b00001000110010: pixel[2:0] = 3'b000;
      14'b00001000110011: pixel[2:0] = 3'b000;
      14'b00001000110100: pixel[2:0] = 3'b000;
      14'b00001000110101: pixel[2:0] = 3'b000;
      14'b00001000110110: pixel[2:0] = 3'b111;
      14'b00001000110111: pixel[2:0] = 3'b111;
      14'b00001000111000: pixel[2:0] = 3'b111;
      14'b00001000111001: pixel[2:0] = 3'b111;
      14'b00001000111010: pixel[2:0] = 3'b000;
      14'b00001000111011: pixel[2:0] = 3'b000;
      14'b00001000111100: pixel[2:0] = 3'b000;
      14'b00001000111101: pixel[2:0] = 3'b000;
      14'b00001000111110: pixel[2:0] = 3'b000;
      14'b00001000111111: pixel[2:0] = 3'b000;
      14'b00001001000000: pixel[2:0] = 3'b000;
      14'b00001001000001: pixel[2:0] = 3'b111;
      14'b00001001000010: pixel[2:0] = 3'b111;
      14'b00001001000011: pixel[2:0] = 3'b111;
      14'b00001001000100: pixel[2:0] = 3'b111;
      14'b00001001000101: pixel[2:0] = 3'b111;
      14'b00001001000110: pixel[2:0] = 3'b000;
      14'b00001001000111: pixel[2:0] = 3'b000;
      14'b00001001001000: pixel[2:0] = 3'b000;
      14'b00001001001001: pixel[2:0] = 3'b000;
      14'b00001001001010: pixel[2:0] = 3'b000;
      14'b00001001001011: pixel[2:0] = 3'b000;
      14'b00001001001100: pixel[2:0] = 3'b000;
      14'b00001001001101: pixel[2:0] = 3'b000;
      14'b00001001001110: pixel[2:0] = 3'b000;
      14'b00001001001111: pixel[2:0] = 3'b000;
      14'b00001001010000: pixel[2:0] = 3'b111;
      14'b00001001010001: pixel[2:0] = 3'b111;
      14'b00001001010010: pixel[2:0] = 3'b111;
      14'b00001001010011: pixel[2:0] = 3'b111;
      14'b00001001010100: pixel[2:0] = 3'b111;
      14'b00001001010101: pixel[2:0] = 3'b111;
      14'b00001001010110: pixel[2:0] = 3'b000;
      14'b00001001010111: pixel[2:0] = 3'b000;
      14'b00001001011000: pixel[2:0] = 3'b000;
      14'b00001001011001: pixel[2:0] = 3'b000;
      14'b00001001011010: pixel[2:0] = 3'b111;
      14'b00001001011011: pixel[2:0] = 3'b111;
      14'b00001001011100: pixel[2:0] = 3'b111;
      14'b00001001011101: pixel[2:0] = 3'b111;
      14'b00001001011110: pixel[2:0] = 3'b111;
      14'b00001001011111: pixel[2:0] = 3'b111;
      14'b00001001100000: pixel[2:0] = 3'b111;
      14'b00001001100001: pixel[2:0] = 3'b111;
      14'b00001001100010: pixel[2:0] = 3'b111;
      14'b00001001100011: pixel[2:0] = 3'b111;
      14'b00001001100100: pixel[2:0] = 3'b111;
      14'b00001001100101: pixel[2:0] = 3'b111;
      14'b00001001100110: pixel[2:0] = 3'b111;
      14'b00001001100111: pixel[2:0] = 3'b111;
      14'b00001001101000: pixel[2:0] = 3'b111;
      14'b00001001101001: pixel[2:0] = 3'b111;
      14'b00001001101010: pixel[2:0] = 3'b111;
      14'b00001001101011: pixel[2:0] = 3'b000;
      14'b00001001101100: pixel[2:0] = 3'b000;
      14'b00001001101101: pixel[2:0] = 3'b000;
      14'b00001001101110: pixel[2:0] = 3'b000;
      14'b00001001101111: pixel[2:0] = 3'b000;
      14'b00001001110000: pixel[2:0] = 3'b111;
      14'b00001001110001: pixel[2:0] = 3'b111;
      14'b00001001110010: pixel[2:0] = 3'b111;
      14'b00001001110011: pixel[2:0] = 3'b111;
      14'b00001001110100: pixel[2:0] = 3'b111;
      14'b00001001110101: pixel[2:0] = 3'b111;
      14'b00001001110110: pixel[2:0] = 3'b111;
      14'b00001001110111: pixel[2:0] = 3'b111;
      14'b00001001111000: pixel[2:0] = 3'b111;
      14'b00001001111001: pixel[2:0] = 3'b111;
      14'b00001001111010: pixel[2:0] = 3'b111;
      14'b00001001111011: pixel[2:0] = 3'b111;
      14'b00001001111100: pixel[2:0] = 3'b000;
      14'b00001001111101: pixel[2:0] = 3'b000;
      14'b00001001111110: pixel[2:0] = 3'b000;
      14'b00001001111111: pixel[2:0] = 3'b000;
      14'b00001010000000: pixel[2:0] = 3'b000;
      14'b00001010000001: pixel[2:0] = 3'b000;
      14'b00001010000010: pixel[2:0] = 3'b000;
      14'b00001010000011: pixel[2:0] = 3'b000;
      14'b00001010000100: pixel[2:0] = 3'b000;
      14'b00001010000101: pixel[2:0] = 3'b000;
      14'b00001010000110: pixel[2:0] = 3'b000;
      14'b00001010000111: pixel[2:0] = 3'b000;
      14'b00001100000000: pixel[2:0] = 3'b000;
      14'b00001100000001: pixel[2:0] = 3'b000;
      14'b00001100000010: pixel[2:0] = 3'b111;
      14'b00001100000011: pixel[2:0] = 3'b111;
      14'b00001100000100: pixel[2:0] = 3'b111;
      14'b00001100000101: pixel[2:0] = 3'b111;
      14'b00001100000110: pixel[2:0] = 3'b111;
      14'b00001100000111: pixel[2:0] = 3'b111;
      14'b00001100001000: pixel[2:0] = 3'b111;
      14'b00001100001001: pixel[2:0] = 3'b111;
      14'b00001100001010: pixel[2:0] = 3'b111;
      14'b00001100001011: pixel[2:0] = 3'b111;
      14'b00001100001100: pixel[2:0] = 3'b111;
      14'b00001100001101: pixel[2:0] = 3'b111;
      14'b00001100001110: pixel[2:0] = 3'b111;
      14'b00001100001111: pixel[2:0] = 3'b111;
      14'b00001100010000: pixel[2:0] = 3'b000;
      14'b00001100010001: pixel[2:0] = 3'b000;
      14'b00001100010010: pixel[2:0] = 3'b000;
      14'b00001100010011: pixel[2:0] = 3'b000;
      14'b00001100010100: pixel[2:0] = 3'b000;
      14'b00001100010101: pixel[2:0] = 3'b000;
      14'b00001100010110: pixel[2:0] = 3'b000;
      14'b00001100010111: pixel[2:0] = 3'b000;
      14'b00001100011000: pixel[2:0] = 3'b000;
      14'b00001100011001: pixel[2:0] = 3'b111;
      14'b00001100011010: pixel[2:0] = 3'b111;
      14'b00001100011011: pixel[2:0] = 3'b111;
      14'b00001100011100: pixel[2:0] = 3'b111;
      14'b00001100011101: pixel[2:0] = 3'b111;
      14'b00001100011110: pixel[2:0] = 3'b000;
      14'b00001100011111: pixel[2:0] = 3'b000;
      14'b00001100100000: pixel[2:0] = 3'b000;
      14'b00001100100001: pixel[2:0] = 3'b000;
      14'b00001100100010: pixel[2:0] = 3'b000;
      14'b00001100100011: pixel[2:0] = 3'b000;
      14'b00001100100100: pixel[2:0] = 3'b000;
      14'b00001100100101: pixel[2:0] = 3'b000;
      14'b00001100100110: pixel[2:0] = 3'b000;
      14'b00001100100111: pixel[2:0] = 3'b000;
      14'b00001100101000: pixel[2:0] = 3'b000;
      14'b00001100101001: pixel[2:0] = 3'b000;
      14'b00001100101010: pixel[2:0] = 3'b000;
      14'b00001100101011: pixel[2:0] = 3'b000;
      14'b00001100101100: pixel[2:0] = 3'b000;
      14'b00001100101101: pixel[2:0] = 3'b000;
      14'b00001100101110: pixel[2:0] = 3'b000;
      14'b00001100101111: pixel[2:0] = 3'b000;
      14'b00001100110000: pixel[2:0] = 3'b000;
      14'b00001100110001: pixel[2:0] = 3'b000;
      14'b00001100110010: pixel[2:0] = 3'b000;
      14'b00001100110011: pixel[2:0] = 3'b000;
      14'b00001100110100: pixel[2:0] = 3'b000;
      14'b00001100110101: pixel[2:0] = 3'b111;
      14'b00001100110110: pixel[2:0] = 3'b111;
      14'b00001100110111: pixel[2:0] = 3'b111;
      14'b00001100111000: pixel[2:0] = 3'b111;
      14'b00001100111001: pixel[2:0] = 3'b111;
      14'b00001100111010: pixel[2:0] = 3'b000;
      14'b00001100111011: pixel[2:0] = 3'b000;
      14'b00001100111100: pixel[2:0] = 3'b000;
      14'b00001100111101: pixel[2:0] = 3'b000;
      14'b00001100111110: pixel[2:0] = 3'b000;
      14'b00001100111111: pixel[2:0] = 3'b000;
      14'b00001101000000: pixel[2:0] = 3'b000;
      14'b00001101000001: pixel[2:0] = 3'b111;
      14'b00001101000010: pixel[2:0] = 3'b111;
      14'b00001101000011: pixel[2:0] = 3'b111;
      14'b00001101000100: pixel[2:0] = 3'b111;
      14'b00001101000101: pixel[2:0] = 3'b111;
      14'b00001101000110: pixel[2:0] = 3'b000;
      14'b00001101000111: pixel[2:0] = 3'b000;
      14'b00001101001000: pixel[2:0] = 3'b000;
      14'b00001101001001: pixel[2:0] = 3'b000;
      14'b00001101001010: pixel[2:0] = 3'b000;
      14'b00001101001011: pixel[2:0] = 3'b000;
      14'b00001101001100: pixel[2:0] = 3'b000;
      14'b00001101001101: pixel[2:0] = 3'b000;
      14'b00001101001110: pixel[2:0] = 3'b000;
      14'b00001101001111: pixel[2:0] = 3'b000;
      14'b00001101010000: pixel[2:0] = 3'b111;
      14'b00001101010001: pixel[2:0] = 3'b111;
      14'b00001101010010: pixel[2:0] = 3'b111;
      14'b00001101010011: pixel[2:0] = 3'b111;
      14'b00001101010100: pixel[2:0] = 3'b111;
      14'b00001101010101: pixel[2:0] = 3'b000;
      14'b00001101010110: pixel[2:0] = 3'b000;
      14'b00001101010111: pixel[2:0] = 3'b000;
      14'b00001101011000: pixel[2:0] = 3'b000;
      14'b00001101011001: pixel[2:0] = 3'b000;
      14'b00001101011010: pixel[2:0] = 3'b111;
      14'b00001101011011: pixel[2:0] = 3'b111;
      14'b00001101011100: pixel[2:0] = 3'b111;
      14'b00001101011101: pixel[2:0] = 3'b111;
      14'b00001101011110: pixel[2:0] = 3'b111;
      14'b00001101011111: pixel[2:0] = 3'b111;
      14'b00001101100000: pixel[2:0] = 3'b111;
      14'b00001101100001: pixel[2:0] = 3'b111;
      14'b00001101100010: pixel[2:0] = 3'b111;
      14'b00001101100011: pixel[2:0] = 3'b111;
      14'b00001101100100: pixel[2:0] = 3'b111;
      14'b00001101100101: pixel[2:0] = 3'b111;
      14'b00001101100110: pixel[2:0] = 3'b111;
      14'b00001101100111: pixel[2:0] = 3'b111;
      14'b00001101101000: pixel[2:0] = 3'b111;
      14'b00001101101001: pixel[2:0] = 3'b111;
      14'b00001101101010: pixel[2:0] = 3'b111;
      14'b00001101101011: pixel[2:0] = 3'b000;
      14'b00001101101100: pixel[2:0] = 3'b000;
      14'b00001101101101: pixel[2:0] = 3'b000;
      14'b00001101101110: pixel[2:0] = 3'b000;
      14'b00001101101111: pixel[2:0] = 3'b000;
      14'b00001101110000: pixel[2:0] = 3'b111;
      14'b00001101110001: pixel[2:0] = 3'b111;
      14'b00001101110010: pixel[2:0] = 3'b111;
      14'b00001101110011: pixel[2:0] = 3'b111;
      14'b00001101110100: pixel[2:0] = 3'b111;
      14'b00001101110101: pixel[2:0] = 3'b111;
      14'b00001101110110: pixel[2:0] = 3'b111;
      14'b00001101110111: pixel[2:0] = 3'b111;
      14'b00001101111000: pixel[2:0] = 3'b111;
      14'b00001101111001: pixel[2:0] = 3'b111;
      14'b00001101111010: pixel[2:0] = 3'b111;
      14'b00001101111011: pixel[2:0] = 3'b111;
      14'b00001101111100: pixel[2:0] = 3'b111;
      14'b00001101111101: pixel[2:0] = 3'b111;
      14'b00001101111110: pixel[2:0] = 3'b000;
      14'b00001101111111: pixel[2:0] = 3'b000;
      14'b00001110000000: pixel[2:0] = 3'b000;
      14'b00001110000001: pixel[2:0] = 3'b000;
      14'b00001110000010: pixel[2:0] = 3'b000;
      14'b00001110000011: pixel[2:0] = 3'b000;
      14'b00001110000100: pixel[2:0] = 3'b000;
      14'b00001110000101: pixel[2:0] = 3'b000;
      14'b00001110000110: pixel[2:0] = 3'b000;
      14'b00001110000111: pixel[2:0] = 3'b000;
      14'b00010000000000: pixel[2:0] = 3'b000;
      14'b00010000000001: pixel[2:0] = 3'b000;
      14'b00010000000010: pixel[2:0] = 3'b111;
      14'b00010000000011: pixel[2:0] = 3'b111;
      14'b00010000000100: pixel[2:0] = 3'b111;
      14'b00010000000101: pixel[2:0] = 3'b111;
      14'b00010000000110: pixel[2:0] = 3'b111;
      14'b00010000000111: pixel[2:0] = 3'b111;
      14'b00010000001000: pixel[2:0] = 3'b111;
      14'b00010000001001: pixel[2:0] = 3'b111;
      14'b00010000001010: pixel[2:0] = 3'b111;
      14'b00010000001011: pixel[2:0] = 3'b111;
      14'b00010000001100: pixel[2:0] = 3'b111;
      14'b00010000001101: pixel[2:0] = 3'b111;
      14'b00010000001110: pixel[2:0] = 3'b111;
      14'b00010000001111: pixel[2:0] = 3'b111;
      14'b00010000010000: pixel[2:0] = 3'b111;
      14'b00010000010001: pixel[2:0] = 3'b000;
      14'b00010000010010: pixel[2:0] = 3'b000;
      14'b00010000010011: pixel[2:0] = 3'b000;
      14'b00010000010100: pixel[2:0] = 3'b000;
      14'b00010000010101: pixel[2:0] = 3'b000;
      14'b00010000010110: pixel[2:0] = 3'b000;
      14'b00010000010111: pixel[2:0] = 3'b000;
      14'b00010000011000: pixel[2:0] = 3'b000;
      14'b00010000011001: pixel[2:0] = 3'b111;
      14'b00010000011010: pixel[2:0] = 3'b111;
      14'b00010000011011: pixel[2:0] = 3'b111;
      14'b00010000011100: pixel[2:0] = 3'b111;
      14'b00010000011101: pixel[2:0] = 3'b111;
      14'b00010000011110: pixel[2:0] = 3'b000;
      14'b00010000011111: pixel[2:0] = 3'b000;
      14'b00010000100000: pixel[2:0] = 3'b000;
      14'b00010000100001: pixel[2:0] = 3'b000;
      14'b00010000100010: pixel[2:0] = 3'b000;
      14'b00010000100011: pixel[2:0] = 3'b000;
      14'b00010000100100: pixel[2:0] = 3'b000;
      14'b00010000100101: pixel[2:0] = 3'b000;
      14'b00010000100110: pixel[2:0] = 3'b000;
      14'b00010000100111: pixel[2:0] = 3'b000;
      14'b00010000101000: pixel[2:0] = 3'b000;
      14'b00010000101001: pixel[2:0] = 3'b000;
      14'b00010000101010: pixel[2:0] = 3'b000;
      14'b00010000101011: pixel[2:0] = 3'b000;
      14'b00010000101100: pixel[2:0] = 3'b000;
      14'b00010000101101: pixel[2:0] = 3'b000;
      14'b00010000101110: pixel[2:0] = 3'b000;
      14'b00010000101111: pixel[2:0] = 3'b000;
      14'b00010000110000: pixel[2:0] = 3'b000;
      14'b00010000110001: pixel[2:0] = 3'b000;
      14'b00010000110010: pixel[2:0] = 3'b000;
      14'b00010000110011: pixel[2:0] = 3'b000;
      14'b00010000110100: pixel[2:0] = 3'b000;
      14'b00010000110101: pixel[2:0] = 3'b111;
      14'b00010000110110: pixel[2:0] = 3'b111;
      14'b00010000110111: pixel[2:0] = 3'b111;
      14'b00010000111000: pixel[2:0] = 3'b111;
      14'b00010000111001: pixel[2:0] = 3'b111;
      14'b00010000111010: pixel[2:0] = 3'b000;
      14'b00010000111011: pixel[2:0] = 3'b000;
      14'b00010000111100: pixel[2:0] = 3'b000;
      14'b00010000111101: pixel[2:0] = 3'b000;
      14'b00010000111110: pixel[2:0] = 3'b000;
      14'b00010000111111: pixel[2:0] = 3'b000;
      14'b00010001000000: pixel[2:0] = 3'b000;
      14'b00010001000001: pixel[2:0] = 3'b000;
      14'b00010001000010: pixel[2:0] = 3'b111;
      14'b00010001000011: pixel[2:0] = 3'b111;
      14'b00010001000100: pixel[2:0] = 3'b111;
      14'b00010001000101: pixel[2:0] = 3'b111;
      14'b00010001000110: pixel[2:0] = 3'b111;
      14'b00010001000111: pixel[2:0] = 3'b000;
      14'b00010001001000: pixel[2:0] = 3'b000;
      14'b00010001001001: pixel[2:0] = 3'b000;
      14'b00010001001010: pixel[2:0] = 3'b000;
      14'b00010001001011: pixel[2:0] = 3'b000;
      14'b00010001001100: pixel[2:0] = 3'b000;
      14'b00010001001101: pixel[2:0] = 3'b000;
      14'b00010001001110: pixel[2:0] = 3'b000;
      14'b00010001001111: pixel[2:0] = 3'b000;
      14'b00010001010000: pixel[2:0] = 3'b111;
      14'b00010001010001: pixel[2:0] = 3'b111;
      14'b00010001010010: pixel[2:0] = 3'b111;
      14'b00010001010011: pixel[2:0] = 3'b111;
      14'b00010001010100: pixel[2:0] = 3'b111;
      14'b00010001010101: pixel[2:0] = 3'b000;
      14'b00010001010110: pixel[2:0] = 3'b000;
      14'b00010001010111: pixel[2:0] = 3'b000;
      14'b00010001011000: pixel[2:0] = 3'b000;
      14'b00010001011001: pixel[2:0] = 3'b000;
      14'b00010001011010: pixel[2:0] = 3'b111;
      14'b00010001011011: pixel[2:0] = 3'b111;
      14'b00010001011100: pixel[2:0] = 3'b111;
      14'b00010001011101: pixel[2:0] = 3'b111;
      14'b00010001011110: pixel[2:0] = 3'b111;
      14'b00010001011111: pixel[2:0] = 3'b111;
      14'b00010001100000: pixel[2:0] = 3'b111;
      14'b00010001100001: pixel[2:0] = 3'b111;
      14'b00010001100010: pixel[2:0] = 3'b111;
      14'b00010001100011: pixel[2:0] = 3'b111;
      14'b00010001100100: pixel[2:0] = 3'b111;
      14'b00010001100101: pixel[2:0] = 3'b111;
      14'b00010001100110: pixel[2:0] = 3'b111;
      14'b00010001100111: pixel[2:0] = 3'b111;
      14'b00010001101000: pixel[2:0] = 3'b111;
      14'b00010001101001: pixel[2:0] = 3'b111;
      14'b00010001101010: pixel[2:0] = 3'b111;
      14'b00010001101011: pixel[2:0] = 3'b000;
      14'b00010001101100: pixel[2:0] = 3'b000;
      14'b00010001101101: pixel[2:0] = 3'b000;
      14'b00010001101110: pixel[2:0] = 3'b000;
      14'b00010001101111: pixel[2:0] = 3'b000;
      14'b00010001110000: pixel[2:0] = 3'b111;
      14'b00010001110001: pixel[2:0] = 3'b111;
      14'b00010001110010: pixel[2:0] = 3'b111;
      14'b00010001110011: pixel[2:0] = 3'b111;
      14'b00010001110100: pixel[2:0] = 3'b111;
      14'b00010001110101: pixel[2:0] = 3'b111;
      14'b00010001110110: pixel[2:0] = 3'b111;
      14'b00010001110111: pixel[2:0] = 3'b111;
      14'b00010001111000: pixel[2:0] = 3'b111;
      14'b00010001111001: pixel[2:0] = 3'b111;
      14'b00010001111010: pixel[2:0] = 3'b111;
      14'b00010001111011: pixel[2:0] = 3'b111;
      14'b00010001111100: pixel[2:0] = 3'b111;
      14'b00010001111101: pixel[2:0] = 3'b111;
      14'b00010001111110: pixel[2:0] = 3'b111;
      14'b00010001111111: pixel[2:0] = 3'b111;
      14'b00010010000000: pixel[2:0] = 3'b000;
      14'b00010010000001: pixel[2:0] = 3'b000;
      14'b00010010000010: pixel[2:0] = 3'b000;
      14'b00010010000011: pixel[2:0] = 3'b000;
      14'b00010010000100: pixel[2:0] = 3'b000;
      14'b00010010000101: pixel[2:0] = 3'b000;
      14'b00010010000110: pixel[2:0] = 3'b000;
      14'b00010010000111: pixel[2:0] = 3'b000;
      14'b00010100000000: pixel[2:0] = 3'b000;
      14'b00010100000001: pixel[2:0] = 3'b000;
      14'b00010100000010: pixel[2:0] = 3'b111;
      14'b00010100000011: pixel[2:0] = 3'b111;
      14'b00010100000100: pixel[2:0] = 3'b111;
      14'b00010100000101: pixel[2:0] = 3'b111;
      14'b00010100000110: pixel[2:0] = 3'b111;
      14'b00010100000111: pixel[2:0] = 3'b111;
      14'b00010100001000: pixel[2:0] = 3'b111;
      14'b00010100001001: pixel[2:0] = 3'b111;
      14'b00010100001010: pixel[2:0] = 3'b111;
      14'b00010100001011: pixel[2:0] = 3'b111;
      14'b00010100001100: pixel[2:0] = 3'b111;
      14'b00010100001101: pixel[2:0] = 3'b111;
      14'b00010100001110: pixel[2:0] = 3'b111;
      14'b00010100001111: pixel[2:0] = 3'b111;
      14'b00010100010000: pixel[2:0] = 3'b111;
      14'b00010100010001: pixel[2:0] = 3'b111;
      14'b00010100010010: pixel[2:0] = 3'b000;
      14'b00010100010011: pixel[2:0] = 3'b000;
      14'b00010100010100: pixel[2:0] = 3'b000;
      14'b00010100010101: pixel[2:0] = 3'b000;
      14'b00010100010110: pixel[2:0] = 3'b000;
      14'b00010100010111: pixel[2:0] = 3'b000;
      14'b00010100011000: pixel[2:0] = 3'b000;
      14'b00010100011001: pixel[2:0] = 3'b111;
      14'b00010100011010: pixel[2:0] = 3'b111;
      14'b00010100011011: pixel[2:0] = 3'b111;
      14'b00010100011100: pixel[2:0] = 3'b111;
      14'b00010100011101: pixel[2:0] = 3'b111;
      14'b00010100011110: pixel[2:0] = 3'b000;
      14'b00010100011111: pixel[2:0] = 3'b000;
      14'b00010100100000: pixel[2:0] = 3'b000;
      14'b00010100100001: pixel[2:0] = 3'b000;
      14'b00010100100010: pixel[2:0] = 3'b000;
      14'b00010100100011: pixel[2:0] = 3'b000;
      14'b00010100100100: pixel[2:0] = 3'b000;
      14'b00010100100101: pixel[2:0] = 3'b000;
      14'b00010100100110: pixel[2:0] = 3'b000;
      14'b00010100100111: pixel[2:0] = 3'b000;
      14'b00010100101000: pixel[2:0] = 3'b000;
      14'b00010100101001: pixel[2:0] = 3'b000;
      14'b00010100101010: pixel[2:0] = 3'b000;
      14'b00010100101011: pixel[2:0] = 3'b000;
      14'b00010100101100: pixel[2:0] = 3'b000;
      14'b00010100101101: pixel[2:0] = 3'b000;
      14'b00010100101110: pixel[2:0] = 3'b000;
      14'b00010100101111: pixel[2:0] = 3'b000;
      14'b00010100110000: pixel[2:0] = 3'b000;
      14'b00010100110001: pixel[2:0] = 3'b000;
      14'b00010100110010: pixel[2:0] = 3'b000;
      14'b00010100110011: pixel[2:0] = 3'b000;
      14'b00010100110100: pixel[2:0] = 3'b000;
      14'b00010100110101: pixel[2:0] = 3'b111;
      14'b00010100110110: pixel[2:0] = 3'b111;
      14'b00010100110111: pixel[2:0] = 3'b111;
      14'b00010100111000: pixel[2:0] = 3'b111;
      14'b00010100111001: pixel[2:0] = 3'b111;
      14'b00010100111010: pixel[2:0] = 3'b111;
      14'b00010100111011: pixel[2:0] = 3'b000;
      14'b00010100111100: pixel[2:0] = 3'b000;
      14'b00010100111101: pixel[2:0] = 3'b000;
      14'b00010100111110: pixel[2:0] = 3'b000;
      14'b00010100111111: pixel[2:0] = 3'b000;
      14'b00010101000000: pixel[2:0] = 3'b000;
      14'b00010101000001: pixel[2:0] = 3'b000;
      14'b00010101000010: pixel[2:0] = 3'b111;
      14'b00010101000011: pixel[2:0] = 3'b111;
      14'b00010101000100: pixel[2:0] = 3'b111;
      14'b00010101000101: pixel[2:0] = 3'b111;
      14'b00010101000110: pixel[2:0] = 3'b111;
      14'b00010101000111: pixel[2:0] = 3'b000;
      14'b00010101001000: pixel[2:0] = 3'b000;
      14'b00010101001001: pixel[2:0] = 3'b000;
      14'b00010101001010: pixel[2:0] = 3'b000;
      14'b00010101001011: pixel[2:0] = 3'b000;
      14'b00010101001100: pixel[2:0] = 3'b000;
      14'b00010101001101: pixel[2:0] = 3'b000;
      14'b00010101001110: pixel[2:0] = 3'b000;
      14'b00010101001111: pixel[2:0] = 3'b000;
      14'b00010101010000: pixel[2:0] = 3'b111;
      14'b00010101010001: pixel[2:0] = 3'b111;
      14'b00010101010010: pixel[2:0] = 3'b111;
      14'b00010101010011: pixel[2:0] = 3'b111;
      14'b00010101010100: pixel[2:0] = 3'b111;
      14'b00010101010101: pixel[2:0] = 3'b000;
      14'b00010101010110: pixel[2:0] = 3'b000;
      14'b00010101010111: pixel[2:0] = 3'b000;
      14'b00010101011000: pixel[2:0] = 3'b000;
      14'b00010101011001: pixel[2:0] = 3'b000;
      14'b00010101011010: pixel[2:0] = 3'b111;
      14'b00010101011011: pixel[2:0] = 3'b111;
      14'b00010101011100: pixel[2:0] = 3'b111;
      14'b00010101011101: pixel[2:0] = 3'b111;
      14'b00010101011110: pixel[2:0] = 3'b111;
      14'b00010101011111: pixel[2:0] = 3'b111;
      14'b00010101100000: pixel[2:0] = 3'b111;
      14'b00010101100001: pixel[2:0] = 3'b111;
      14'b00010101100010: pixel[2:0] = 3'b111;
      14'b00010101100011: pixel[2:0] = 3'b111;
      14'b00010101100100: pixel[2:0] = 3'b111;
      14'b00010101100101: pixel[2:0] = 3'b111;
      14'b00010101100110: pixel[2:0] = 3'b111;
      14'b00010101100111: pixel[2:0] = 3'b111;
      14'b00010101101000: pixel[2:0] = 3'b111;
      14'b00010101101001: pixel[2:0] = 3'b111;
      14'b00010101101010: pixel[2:0] = 3'b111;
      14'b00010101101011: pixel[2:0] = 3'b000;
      14'b00010101101100: pixel[2:0] = 3'b000;
      14'b00010101101101: pixel[2:0] = 3'b000;
      14'b00010101101110: pixel[2:0] = 3'b000;
      14'b00010101101111: pixel[2:0] = 3'b000;
      14'b00010101110000: pixel[2:0] = 3'b111;
      14'b00010101110001: pixel[2:0] = 3'b111;
      14'b00010101110010: pixel[2:0] = 3'b111;
      14'b00010101110011: pixel[2:0] = 3'b111;
      14'b00010101110100: pixel[2:0] = 3'b111;
      14'b00010101110101: pixel[2:0] = 3'b111;
      14'b00010101110110: pixel[2:0] = 3'b111;
      14'b00010101110111: pixel[2:0] = 3'b111;
      14'b00010101111000: pixel[2:0] = 3'b111;
      14'b00010101111001: pixel[2:0] = 3'b111;
      14'b00010101111010: pixel[2:0] = 3'b111;
      14'b00010101111011: pixel[2:0] = 3'b111;
      14'b00010101111100: pixel[2:0] = 3'b111;
      14'b00010101111101: pixel[2:0] = 3'b111;
      14'b00010101111110: pixel[2:0] = 3'b111;
      14'b00010101111111: pixel[2:0] = 3'b111;
      14'b00010110000000: pixel[2:0] = 3'b111;
      14'b00010110000001: pixel[2:0] = 3'b000;
      14'b00010110000010: pixel[2:0] = 3'b000;
      14'b00010110000011: pixel[2:0] = 3'b000;
      14'b00010110000100: pixel[2:0] = 3'b000;
      14'b00010110000101: pixel[2:0] = 3'b000;
      14'b00010110000110: pixel[2:0] = 3'b000;
      14'b00010110000111: pixel[2:0] = 3'b000;
      14'b00011000000000: pixel[2:0] = 3'b000;
      14'b00011000000001: pixel[2:0] = 3'b000;
      14'b00011000000010: pixel[2:0] = 3'b111;
      14'b00011000000011: pixel[2:0] = 3'b111;
      14'b00011000000100: pixel[2:0] = 3'b111;
      14'b00011000000101: pixel[2:0] = 3'b111;
      14'b00011000000110: pixel[2:0] = 3'b111;
      14'b00011000000111: pixel[2:0] = 3'b111;
      14'b00011000001000: pixel[2:0] = 3'b111;
      14'b00011000001001: pixel[2:0] = 3'b111;
      14'b00011000001010: pixel[2:0] = 3'b111;
      14'b00011000001011: pixel[2:0] = 3'b111;
      14'b00011000001100: pixel[2:0] = 3'b111;
      14'b00011000001101: pixel[2:0] = 3'b111;
      14'b00011000001110: pixel[2:0] = 3'b111;
      14'b00011000001111: pixel[2:0] = 3'b111;
      14'b00011000010000: pixel[2:0] = 3'b111;
      14'b00011000010001: pixel[2:0] = 3'b111;
      14'b00011000010010: pixel[2:0] = 3'b111;
      14'b00011000010011: pixel[2:0] = 3'b000;
      14'b00011000010100: pixel[2:0] = 3'b000;
      14'b00011000010101: pixel[2:0] = 3'b000;
      14'b00011000010110: pixel[2:0] = 3'b000;
      14'b00011000010111: pixel[2:0] = 3'b000;
      14'b00011000011000: pixel[2:0] = 3'b000;
      14'b00011000011001: pixel[2:0] = 3'b111;
      14'b00011000011010: pixel[2:0] = 3'b111;
      14'b00011000011011: pixel[2:0] = 3'b111;
      14'b00011000011100: pixel[2:0] = 3'b111;
      14'b00011000011101: pixel[2:0] = 3'b111;
      14'b00011000011110: pixel[2:0] = 3'b000;
      14'b00011000011111: pixel[2:0] = 3'b000;
      14'b00011000100000: pixel[2:0] = 3'b000;
      14'b00011000100001: pixel[2:0] = 3'b000;
      14'b00011000100010: pixel[2:0] = 3'b000;
      14'b00011000100011: pixel[2:0] = 3'b000;
      14'b00011000100100: pixel[2:0] = 3'b000;
      14'b00011000100101: pixel[2:0] = 3'b000;
      14'b00011000100110: pixel[2:0] = 3'b000;
      14'b00011000100111: pixel[2:0] = 3'b000;
      14'b00011000101000: pixel[2:0] = 3'b000;
      14'b00011000101001: pixel[2:0] = 3'b000;
      14'b00011000101010: pixel[2:0] = 3'b000;
      14'b00011000101011: pixel[2:0] = 3'b000;
      14'b00011000101100: pixel[2:0] = 3'b000;
      14'b00011000101101: pixel[2:0] = 3'b000;
      14'b00011000101110: pixel[2:0] = 3'b000;
      14'b00011000101111: pixel[2:0] = 3'b000;
      14'b00011000110000: pixel[2:0] = 3'b000;
      14'b00011000110001: pixel[2:0] = 3'b000;
      14'b00011000110010: pixel[2:0] = 3'b000;
      14'b00011000110011: pixel[2:0] = 3'b000;
      14'b00011000110100: pixel[2:0] = 3'b000;
      14'b00011000110101: pixel[2:0] = 3'b111;
      14'b00011000110110: pixel[2:0] = 3'b111;
      14'b00011000110111: pixel[2:0] = 3'b111;
      14'b00011000111000: pixel[2:0] = 3'b111;
      14'b00011000111001: pixel[2:0] = 3'b111;
      14'b00011000111010: pixel[2:0] = 3'b111;
      14'b00011000111011: pixel[2:0] = 3'b000;
      14'b00011000111100: pixel[2:0] = 3'b000;
      14'b00011000111101: pixel[2:0] = 3'b000;
      14'b00011000111110: pixel[2:0] = 3'b000;
      14'b00011000111111: pixel[2:0] = 3'b000;
      14'b00011001000000: pixel[2:0] = 3'b000;
      14'b00011001000001: pixel[2:0] = 3'b000;
      14'b00011001000010: pixel[2:0] = 3'b111;
      14'b00011001000011: pixel[2:0] = 3'b111;
      14'b00011001000100: pixel[2:0] = 3'b111;
      14'b00011001000101: pixel[2:0] = 3'b111;
      14'b00011001000110: pixel[2:0] = 3'b111;
      14'b00011001000111: pixel[2:0] = 3'b000;
      14'b00011001001000: pixel[2:0] = 3'b000;
      14'b00011001001001: pixel[2:0] = 3'b000;
      14'b00011001001010: pixel[2:0] = 3'b000;
      14'b00011001001011: pixel[2:0] = 3'b000;
      14'b00011001001100: pixel[2:0] = 3'b000;
      14'b00011001001101: pixel[2:0] = 3'b000;
      14'b00011001001110: pixel[2:0] = 3'b000;
      14'b00011001001111: pixel[2:0] = 3'b111;
      14'b00011001010000: pixel[2:0] = 3'b111;
      14'b00011001010001: pixel[2:0] = 3'b111;
      14'b00011001010010: pixel[2:0] = 3'b111;
      14'b00011001010011: pixel[2:0] = 3'b111;
      14'b00011001010100: pixel[2:0] = 3'b000;
      14'b00011001010101: pixel[2:0] = 3'b000;
      14'b00011001010110: pixel[2:0] = 3'b000;
      14'b00011001010111: pixel[2:0] = 3'b000;
      14'b00011001011000: pixel[2:0] = 3'b000;
      14'b00011001011001: pixel[2:0] = 3'b000;
      14'b00011001011010: pixel[2:0] = 3'b111;
      14'b00011001011011: pixel[2:0] = 3'b111;
      14'b00011001011100: pixel[2:0] = 3'b111;
      14'b00011001011101: pixel[2:0] = 3'b111;
      14'b00011001011110: pixel[2:0] = 3'b111;
      14'b00011001011111: pixel[2:0] = 3'b111;
      14'b00011001100000: pixel[2:0] = 3'b111;
      14'b00011001100001: pixel[2:0] = 3'b111;
      14'b00011001100010: pixel[2:0] = 3'b111;
      14'b00011001100011: pixel[2:0] = 3'b111;
      14'b00011001100100: pixel[2:0] = 3'b111;
      14'b00011001100101: pixel[2:0] = 3'b111;
      14'b00011001100110: pixel[2:0] = 3'b111;
      14'b00011001100111: pixel[2:0] = 3'b111;
      14'b00011001101000: pixel[2:0] = 3'b111;
      14'b00011001101001: pixel[2:0] = 3'b111;
      14'b00011001101010: pixel[2:0] = 3'b111;
      14'b00011001101011: pixel[2:0] = 3'b000;
      14'b00011001101100: pixel[2:0] = 3'b000;
      14'b00011001101101: pixel[2:0] = 3'b000;
      14'b00011001101110: pixel[2:0] = 3'b000;
      14'b00011001101111: pixel[2:0] = 3'b000;
      14'b00011001110000: pixel[2:0] = 3'b111;
      14'b00011001110001: pixel[2:0] = 3'b111;
      14'b00011001110010: pixel[2:0] = 3'b111;
      14'b00011001110011: pixel[2:0] = 3'b111;
      14'b00011001110100: pixel[2:0] = 3'b111;
      14'b00011001110101: pixel[2:0] = 3'b111;
      14'b00011001110110: pixel[2:0] = 3'b111;
      14'b00011001110111: pixel[2:0] = 3'b111;
      14'b00011001111000: pixel[2:0] = 3'b111;
      14'b00011001111001: pixel[2:0] = 3'b111;
      14'b00011001111010: pixel[2:0] = 3'b111;
      14'b00011001111011: pixel[2:0] = 3'b111;
      14'b00011001111100: pixel[2:0] = 3'b111;
      14'b00011001111101: pixel[2:0] = 3'b111;
      14'b00011001111110: pixel[2:0] = 3'b111;
      14'b00011001111111: pixel[2:0] = 3'b111;
      14'b00011010000000: pixel[2:0] = 3'b111;
      14'b00011010000001: pixel[2:0] = 3'b111;
      14'b00011010000010: pixel[2:0] = 3'b000;
      14'b00011010000011: pixel[2:0] = 3'b000;
      14'b00011010000100: pixel[2:0] = 3'b000;
      14'b00011010000101: pixel[2:0] = 3'b000;
      14'b00011010000110: pixel[2:0] = 3'b000;
      14'b00011010000111: pixel[2:0] = 3'b000;
      14'b00011100000000: pixel[2:0] = 3'b000;
      14'b00011100000001: pixel[2:0] = 3'b000;
      14'b00011100000010: pixel[2:0] = 3'b111;
      14'b00011100000011: pixel[2:0] = 3'b111;
      14'b00011100000100: pixel[2:0] = 3'b111;
      14'b00011100000101: pixel[2:0] = 3'b111;
      14'b00011100000110: pixel[2:0] = 3'b111;
      14'b00011100000111: pixel[2:0] = 3'b111;
      14'b00011100001000: pixel[2:0] = 3'b111;
      14'b00011100001001: pixel[2:0] = 3'b111;
      14'b00011100001010: pixel[2:0] = 3'b111;
      14'b00011100001011: pixel[2:0] = 3'b111;
      14'b00011100001100: pixel[2:0] = 3'b111;
      14'b00011100001101: pixel[2:0] = 3'b111;
      14'b00011100001110: pixel[2:0] = 3'b111;
      14'b00011100001111: pixel[2:0] = 3'b111;
      14'b00011100010000: pixel[2:0] = 3'b111;
      14'b00011100010001: pixel[2:0] = 3'b111;
      14'b00011100010010: pixel[2:0] = 3'b111;
      14'b00011100010011: pixel[2:0] = 3'b000;
      14'b00011100010100: pixel[2:0] = 3'b000;
      14'b00011100010101: pixel[2:0] = 3'b000;
      14'b00011100010110: pixel[2:0] = 3'b000;
      14'b00011100010111: pixel[2:0] = 3'b000;
      14'b00011100011000: pixel[2:0] = 3'b000;
      14'b00011100011001: pixel[2:0] = 3'b111;
      14'b00011100011010: pixel[2:0] = 3'b111;
      14'b00011100011011: pixel[2:0] = 3'b111;
      14'b00011100011100: pixel[2:0] = 3'b111;
      14'b00011100011101: pixel[2:0] = 3'b111;
      14'b00011100011110: pixel[2:0] = 3'b000;
      14'b00011100011111: pixel[2:0] = 3'b000;
      14'b00011100100000: pixel[2:0] = 3'b000;
      14'b00011100100001: pixel[2:0] = 3'b000;
      14'b00011100100010: pixel[2:0] = 3'b000;
      14'b00011100100011: pixel[2:0] = 3'b000;
      14'b00011100100100: pixel[2:0] = 3'b000;
      14'b00011100100101: pixel[2:0] = 3'b000;
      14'b00011100100110: pixel[2:0] = 3'b000;
      14'b00011100100111: pixel[2:0] = 3'b000;
      14'b00011100101000: pixel[2:0] = 3'b000;
      14'b00011100101001: pixel[2:0] = 3'b000;
      14'b00011100101010: pixel[2:0] = 3'b000;
      14'b00011100101011: pixel[2:0] = 3'b000;
      14'b00011100101100: pixel[2:0] = 3'b000;
      14'b00011100101101: pixel[2:0] = 3'b000;
      14'b00011100101110: pixel[2:0] = 3'b000;
      14'b00011100101111: pixel[2:0] = 3'b000;
      14'b00011100110000: pixel[2:0] = 3'b000;
      14'b00011100110001: pixel[2:0] = 3'b000;
      14'b00011100110010: pixel[2:0] = 3'b000;
      14'b00011100110011: pixel[2:0] = 3'b000;
      14'b00011100110100: pixel[2:0] = 3'b000;
      14'b00011100110101: pixel[2:0] = 3'b111;
      14'b00011100110110: pixel[2:0] = 3'b111;
      14'b00011100110111: pixel[2:0] = 3'b111;
      14'b00011100111000: pixel[2:0] = 3'b111;
      14'b00011100111001: pixel[2:0] = 3'b111;
      14'b00011100111010: pixel[2:0] = 3'b111;
      14'b00011100111011: pixel[2:0] = 3'b000;
      14'b00011100111100: pixel[2:0] = 3'b000;
      14'b00011100111101: pixel[2:0] = 3'b000;
      14'b00011100111110: pixel[2:0] = 3'b000;
      14'b00011100111111: pixel[2:0] = 3'b000;
      14'b00011101000000: pixel[2:0] = 3'b000;
      14'b00011101000001: pixel[2:0] = 3'b000;
      14'b00011101000010: pixel[2:0] = 3'b000;
      14'b00011101000011: pixel[2:0] = 3'b111;
      14'b00011101000100: pixel[2:0] = 3'b111;
      14'b00011101000101: pixel[2:0] = 3'b111;
      14'b00011101000110: pixel[2:0] = 3'b111;
      14'b00011101000111: pixel[2:0] = 3'b111;
      14'b00011101001000: pixel[2:0] = 3'b000;
      14'b00011101001001: pixel[2:0] = 3'b000;
      14'b00011101001010: pixel[2:0] = 3'b000;
      14'b00011101001011: pixel[2:0] = 3'b000;
      14'b00011101001100: pixel[2:0] = 3'b000;
      14'b00011101001101: pixel[2:0] = 3'b000;
      14'b00011101001110: pixel[2:0] = 3'b000;
      14'b00011101001111: pixel[2:0] = 3'b111;
      14'b00011101010000: pixel[2:0] = 3'b111;
      14'b00011101010001: pixel[2:0] = 3'b111;
      14'b00011101010010: pixel[2:0] = 3'b111;
      14'b00011101010011: pixel[2:0] = 3'b111;
      14'b00011101010100: pixel[2:0] = 3'b000;
      14'b00011101010101: pixel[2:0] = 3'b000;
      14'b00011101010110: pixel[2:0] = 3'b000;
      14'b00011101010111: pixel[2:0] = 3'b000;
      14'b00011101011000: pixel[2:0] = 3'b000;
      14'b00011101011001: pixel[2:0] = 3'b000;
      14'b00011101011010: pixel[2:0] = 3'b111;
      14'b00011101011011: pixel[2:0] = 3'b111;
      14'b00011101011100: pixel[2:0] = 3'b111;
      14'b00011101011101: pixel[2:0] = 3'b111;
      14'b00011101011110: pixel[2:0] = 3'b111;
      14'b00011101011111: pixel[2:0] = 3'b111;
      14'b00011101100000: pixel[2:0] = 3'b111;
      14'b00011101100001: pixel[2:0] = 3'b111;
      14'b00011101100010: pixel[2:0] = 3'b111;
      14'b00011101100011: pixel[2:0] = 3'b111;
      14'b00011101100100: pixel[2:0] = 3'b111;
      14'b00011101100101: pixel[2:0] = 3'b111;
      14'b00011101100110: pixel[2:0] = 3'b111;
      14'b00011101100111: pixel[2:0] = 3'b111;
      14'b00011101101000: pixel[2:0] = 3'b111;
      14'b00011101101001: pixel[2:0] = 3'b111;
      14'b00011101101010: pixel[2:0] = 3'b111;
      14'b00011101101011: pixel[2:0] = 3'b000;
      14'b00011101101100: pixel[2:0] = 3'b000;
      14'b00011101101101: pixel[2:0] = 3'b000;
      14'b00011101101110: pixel[2:0] = 3'b000;
      14'b00011101101111: pixel[2:0] = 3'b000;
      14'b00011101110000: pixel[2:0] = 3'b111;
      14'b00011101110001: pixel[2:0] = 3'b111;
      14'b00011101110010: pixel[2:0] = 3'b111;
      14'b00011101110011: pixel[2:0] = 3'b111;
      14'b00011101110100: pixel[2:0] = 3'b111;
      14'b00011101110101: pixel[2:0] = 3'b111;
      14'b00011101110110: pixel[2:0] = 3'b111;
      14'b00011101110111: pixel[2:0] = 3'b111;
      14'b00011101111000: pixel[2:0] = 3'b111;
      14'b00011101111001: pixel[2:0] = 3'b111;
      14'b00011101111010: pixel[2:0] = 3'b111;
      14'b00011101111011: pixel[2:0] = 3'b111;
      14'b00011101111100: pixel[2:0] = 3'b111;
      14'b00011101111101: pixel[2:0] = 3'b111;
      14'b00011101111110: pixel[2:0] = 3'b111;
      14'b00011101111111: pixel[2:0] = 3'b111;
      14'b00011110000000: pixel[2:0] = 3'b111;
      14'b00011110000001: pixel[2:0] = 3'b111;
      14'b00011110000010: pixel[2:0] = 3'b000;
      14'b00011110000011: pixel[2:0] = 3'b000;
      14'b00011110000100: pixel[2:0] = 3'b000;
      14'b00011110000101: pixel[2:0] = 3'b000;
      14'b00011110000110: pixel[2:0] = 3'b000;
      14'b00011110000111: pixel[2:0] = 3'b000;
      14'b00100000000000: pixel[2:0] = 3'b000;
      14'b00100000000001: pixel[2:0] = 3'b000;
      14'b00100000000010: pixel[2:0] = 3'b111;
      14'b00100000000011: pixel[2:0] = 3'b111;
      14'b00100000000100: pixel[2:0] = 3'b111;
      14'b00100000000101: pixel[2:0] = 3'b111;
      14'b00100000000110: pixel[2:0] = 3'b111;
      14'b00100000000111: pixel[2:0] = 3'b000;
      14'b00100000001000: pixel[2:0] = 3'b000;
      14'b00100000001001: pixel[2:0] = 3'b000;
      14'b00100000001010: pixel[2:0] = 3'b000;
      14'b00100000001011: pixel[2:0] = 3'b000;
      14'b00100000001100: pixel[2:0] = 3'b000;
      14'b00100000001101: pixel[2:0] = 3'b000;
      14'b00100000001110: pixel[2:0] = 3'b111;
      14'b00100000001111: pixel[2:0] = 3'b111;
      14'b00100000010000: pixel[2:0] = 3'b111;
      14'b00100000010001: pixel[2:0] = 3'b111;
      14'b00100000010010: pixel[2:0] = 3'b111;
      14'b00100000010011: pixel[2:0] = 3'b111;
      14'b00100000010100: pixel[2:0] = 3'b000;
      14'b00100000010101: pixel[2:0] = 3'b000;
      14'b00100000010110: pixel[2:0] = 3'b000;
      14'b00100000010111: pixel[2:0] = 3'b000;
      14'b00100000011000: pixel[2:0] = 3'b000;
      14'b00100000011001: pixel[2:0] = 3'b111;
      14'b00100000011010: pixel[2:0] = 3'b111;
      14'b00100000011011: pixel[2:0] = 3'b111;
      14'b00100000011100: pixel[2:0] = 3'b111;
      14'b00100000011101: pixel[2:0] = 3'b111;
      14'b00100000011110: pixel[2:0] = 3'b000;
      14'b00100000011111: pixel[2:0] = 3'b000;
      14'b00100000100000: pixel[2:0] = 3'b000;
      14'b00100000100001: pixel[2:0] = 3'b000;
      14'b00100000100010: pixel[2:0] = 3'b000;
      14'b00100000100011: pixel[2:0] = 3'b000;
      14'b00100000100100: pixel[2:0] = 3'b000;
      14'b00100000100101: pixel[2:0] = 3'b000;
      14'b00100000100110: pixel[2:0] = 3'b000;
      14'b00100000100111: pixel[2:0] = 3'b000;
      14'b00100000101000: pixel[2:0] = 3'b000;
      14'b00100000101001: pixel[2:0] = 3'b000;
      14'b00100000101010: pixel[2:0] = 3'b000;
      14'b00100000101011: pixel[2:0] = 3'b000;
      14'b00100000101100: pixel[2:0] = 3'b000;
      14'b00100000101101: pixel[2:0] = 3'b000;
      14'b00100000101110: pixel[2:0] = 3'b000;
      14'b00100000101111: pixel[2:0] = 3'b000;
      14'b00100000110000: pixel[2:0] = 3'b000;
      14'b00100000110001: pixel[2:0] = 3'b000;
      14'b00100000110010: pixel[2:0] = 3'b000;
      14'b00100000110011: pixel[2:0] = 3'b000;
      14'b00100000110100: pixel[2:0] = 3'b111;
      14'b00100000110101: pixel[2:0] = 3'b111;
      14'b00100000110110: pixel[2:0] = 3'b111;
      14'b00100000110111: pixel[2:0] = 3'b111;
      14'b00100000111000: pixel[2:0] = 3'b111;
      14'b00100000111001: pixel[2:0] = 3'b111;
      14'b00100000111010: pixel[2:0] = 3'b111;
      14'b00100000111011: pixel[2:0] = 3'b000;
      14'b00100000111100: pixel[2:0] = 3'b000;
      14'b00100000111101: pixel[2:0] = 3'b000;
      14'b00100000111110: pixel[2:0] = 3'b000;
      14'b00100000111111: pixel[2:0] = 3'b000;
      14'b00100001000000: pixel[2:0] = 3'b000;
      14'b00100001000001: pixel[2:0] = 3'b000;
      14'b00100001000010: pixel[2:0] = 3'b000;
      14'b00100001000011: pixel[2:0] = 3'b111;
      14'b00100001000100: pixel[2:0] = 3'b111;
      14'b00100001000101: pixel[2:0] = 3'b111;
      14'b00100001000110: pixel[2:0] = 3'b111;
      14'b00100001000111: pixel[2:0] = 3'b111;
      14'b00100001001000: pixel[2:0] = 3'b000;
      14'b00100001001001: pixel[2:0] = 3'b000;
      14'b00100001001010: pixel[2:0] = 3'b000;
      14'b00100001001011: pixel[2:0] = 3'b000;
      14'b00100001001100: pixel[2:0] = 3'b000;
      14'b00100001001101: pixel[2:0] = 3'b000;
      14'b00100001001110: pixel[2:0] = 3'b000;
      14'b00100001001111: pixel[2:0] = 3'b111;
      14'b00100001010000: pixel[2:0] = 3'b111;
      14'b00100001010001: pixel[2:0] = 3'b111;
      14'b00100001010010: pixel[2:0] = 3'b111;
      14'b00100001010011: pixel[2:0] = 3'b111;
      14'b00100001010100: pixel[2:0] = 3'b000;
      14'b00100001010101: pixel[2:0] = 3'b000;
      14'b00100001010110: pixel[2:0] = 3'b000;
      14'b00100001010111: pixel[2:0] = 3'b000;
      14'b00100001011000: pixel[2:0] = 3'b000;
      14'b00100001011001: pixel[2:0] = 3'b000;
      14'b00100001011010: pixel[2:0] = 3'b111;
      14'b00100001011011: pixel[2:0] = 3'b111;
      14'b00100001011100: pixel[2:0] = 3'b111;
      14'b00100001011101: pixel[2:0] = 3'b111;
      14'b00100001011110: pixel[2:0] = 3'b111;
      14'b00100001011111: pixel[2:0] = 3'b000;
      14'b00100001100000: pixel[2:0] = 3'b000;
      14'b00100001100001: pixel[2:0] = 3'b000;
      14'b00100001100010: pixel[2:0] = 3'b000;
      14'b00100001100011: pixel[2:0] = 3'b000;
      14'b00100001100100: pixel[2:0] = 3'b000;
      14'b00100001100101: pixel[2:0] = 3'b000;
      14'b00100001100110: pixel[2:0] = 3'b000;
      14'b00100001100111: pixel[2:0] = 3'b000;
      14'b00100001101000: pixel[2:0] = 3'b000;
      14'b00100001101001: pixel[2:0] = 3'b000;
      14'b00100001101010: pixel[2:0] = 3'b000;
      14'b00100001101011: pixel[2:0] = 3'b000;
      14'b00100001101100: pixel[2:0] = 3'b000;
      14'b00100001101101: pixel[2:0] = 3'b000;
      14'b00100001101110: pixel[2:0] = 3'b000;
      14'b00100001101111: pixel[2:0] = 3'b000;
      14'b00100001110000: pixel[2:0] = 3'b111;
      14'b00100001110001: pixel[2:0] = 3'b111;
      14'b00100001110010: pixel[2:0] = 3'b111;
      14'b00100001110011: pixel[2:0] = 3'b111;
      14'b00100001110100: pixel[2:0] = 3'b111;
      14'b00100001110101: pixel[2:0] = 3'b000;
      14'b00100001110110: pixel[2:0] = 3'b000;
      14'b00100001110111: pixel[2:0] = 3'b000;
      14'b00100001111000: pixel[2:0] = 3'b000;
      14'b00100001111001: pixel[2:0] = 3'b000;
      14'b00100001111010: pixel[2:0] = 3'b000;
      14'b00100001111011: pixel[2:0] = 3'b000;
      14'b00100001111100: pixel[2:0] = 3'b000;
      14'b00100001111101: pixel[2:0] = 3'b111;
      14'b00100001111110: pixel[2:0] = 3'b111;
      14'b00100001111111: pixel[2:0] = 3'b111;
      14'b00100010000000: pixel[2:0] = 3'b111;
      14'b00100010000001: pixel[2:0] = 3'b111;
      14'b00100010000010: pixel[2:0] = 3'b000;
      14'b00100010000011: pixel[2:0] = 3'b000;
      14'b00100010000100: pixel[2:0] = 3'b000;
      14'b00100010000101: pixel[2:0] = 3'b000;
      14'b00100010000110: pixel[2:0] = 3'b000;
      14'b00100010000111: pixel[2:0] = 3'b000;
      14'b00100100000000: pixel[2:0] = 3'b000;
      14'b00100100000001: pixel[2:0] = 3'b000;
      14'b00100100000010: pixel[2:0] = 3'b111;
      14'b00100100000011: pixel[2:0] = 3'b111;
      14'b00100100000100: pixel[2:0] = 3'b111;
      14'b00100100000101: pixel[2:0] = 3'b111;
      14'b00100100000110: pixel[2:0] = 3'b111;
      14'b00100100000111: pixel[2:0] = 3'b000;
      14'b00100100001000: pixel[2:0] = 3'b000;
      14'b00100100001001: pixel[2:0] = 3'b000;
      14'b00100100001010: pixel[2:0] = 3'b000;
      14'b00100100001011: pixel[2:0] = 3'b000;
      14'b00100100001100: pixel[2:0] = 3'b000;
      14'b00100100001101: pixel[2:0] = 3'b000;
      14'b00100100001110: pixel[2:0] = 3'b000;
      14'b00100100001111: pixel[2:0] = 3'b111;
      14'b00100100010000: pixel[2:0] = 3'b111;
      14'b00100100010001: pixel[2:0] = 3'b111;
      14'b00100100010010: pixel[2:0] = 3'b111;
      14'b00100100010011: pixel[2:0] = 3'b111;
      14'b00100100010100: pixel[2:0] = 3'b000;
      14'b00100100010101: pixel[2:0] = 3'b000;
      14'b00100100010110: pixel[2:0] = 3'b000;
      14'b00100100010111: pixel[2:0] = 3'b000;
      14'b00100100011000: pixel[2:0] = 3'b000;
      14'b00100100011001: pixel[2:0] = 3'b111;
      14'b00100100011010: pixel[2:0] = 3'b111;
      14'b00100100011011: pixel[2:0] = 3'b111;
      14'b00100100011100: pixel[2:0] = 3'b111;
      14'b00100100011101: pixel[2:0] = 3'b111;
      14'b00100100011110: pixel[2:0] = 3'b000;
      14'b00100100011111: pixel[2:0] = 3'b000;
      14'b00100100100000: pixel[2:0] = 3'b000;
      14'b00100100100001: pixel[2:0] = 3'b000;
      14'b00100100100010: pixel[2:0] = 3'b000;
      14'b00100100100011: pixel[2:0] = 3'b000;
      14'b00100100100100: pixel[2:0] = 3'b000;
      14'b00100100100101: pixel[2:0] = 3'b000;
      14'b00100100100110: pixel[2:0] = 3'b000;
      14'b00100100100111: pixel[2:0] = 3'b000;
      14'b00100100101000: pixel[2:0] = 3'b000;
      14'b00100100101001: pixel[2:0] = 3'b000;
      14'b00100100101010: pixel[2:0] = 3'b000;
      14'b00100100101011: pixel[2:0] = 3'b000;
      14'b00100100101100: pixel[2:0] = 3'b000;
      14'b00100100101101: pixel[2:0] = 3'b000;
      14'b00100100101110: pixel[2:0] = 3'b000;
      14'b00100100101111: pixel[2:0] = 3'b000;
      14'b00100100110000: pixel[2:0] = 3'b000;
      14'b00100100110001: pixel[2:0] = 3'b000;
      14'b00100100110010: pixel[2:0] = 3'b000;
      14'b00100100110011: pixel[2:0] = 3'b000;
      14'b00100100110100: pixel[2:0] = 3'b111;
      14'b00100100110101: pixel[2:0] = 3'b111;
      14'b00100100110110: pixel[2:0] = 3'b111;
      14'b00100100110111: pixel[2:0] = 3'b111;
      14'b00100100111000: pixel[2:0] = 3'b111;
      14'b00100100111001: pixel[2:0] = 3'b111;
      14'b00100100111010: pixel[2:0] = 3'b111;
      14'b00100100111011: pixel[2:0] = 3'b000;
      14'b00100100111100: pixel[2:0] = 3'b000;
      14'b00100100111101: pixel[2:0] = 3'b000;
      14'b00100100111110: pixel[2:0] = 3'b000;
      14'b00100100111111: pixel[2:0] = 3'b000;
      14'b00100101000000: pixel[2:0] = 3'b000;
      14'b00100101000001: pixel[2:0] = 3'b000;
      14'b00100101000010: pixel[2:0] = 3'b000;
      14'b00100101000011: pixel[2:0] = 3'b111;
      14'b00100101000100: pixel[2:0] = 3'b111;
      14'b00100101000101: pixel[2:0] = 3'b111;
      14'b00100101000110: pixel[2:0] = 3'b111;
      14'b00100101000111: pixel[2:0] = 3'b111;
      14'b00100101001000: pixel[2:0] = 3'b000;
      14'b00100101001001: pixel[2:0] = 3'b000;
      14'b00100101001010: pixel[2:0] = 3'b000;
      14'b00100101001011: pixel[2:0] = 3'b000;
      14'b00100101001100: pixel[2:0] = 3'b000;
      14'b00100101001101: pixel[2:0] = 3'b000;
      14'b00100101001110: pixel[2:0] = 3'b111;
      14'b00100101001111: pixel[2:0] = 3'b111;
      14'b00100101010000: pixel[2:0] = 3'b111;
      14'b00100101010001: pixel[2:0] = 3'b111;
      14'b00100101010010: pixel[2:0] = 3'b111;
      14'b00100101010011: pixel[2:0] = 3'b000;
      14'b00100101010100: pixel[2:0] = 3'b000;
      14'b00100101010101: pixel[2:0] = 3'b000;
      14'b00100101010110: pixel[2:0] = 3'b000;
      14'b00100101010111: pixel[2:0] = 3'b000;
      14'b00100101011000: pixel[2:0] = 3'b000;
      14'b00100101011001: pixel[2:0] = 3'b000;
      14'b00100101011010: pixel[2:0] = 3'b111;
      14'b00100101011011: pixel[2:0] = 3'b111;
      14'b00100101011100: pixel[2:0] = 3'b111;
      14'b00100101011101: pixel[2:0] = 3'b111;
      14'b00100101011110: pixel[2:0] = 3'b111;
      14'b00100101011111: pixel[2:0] = 3'b000;
      14'b00100101100000: pixel[2:0] = 3'b000;
      14'b00100101100001: pixel[2:0] = 3'b000;
      14'b00100101100010: pixel[2:0] = 3'b000;
      14'b00100101100011: pixel[2:0] = 3'b000;
      14'b00100101100100: pixel[2:0] = 3'b000;
      14'b00100101100101: pixel[2:0] = 3'b000;
      14'b00100101100110: pixel[2:0] = 3'b000;
      14'b00100101100111: pixel[2:0] = 3'b000;
      14'b00100101101000: pixel[2:0] = 3'b000;
      14'b00100101101001: pixel[2:0] = 3'b000;
      14'b00100101101010: pixel[2:0] = 3'b000;
      14'b00100101101011: pixel[2:0] = 3'b000;
      14'b00100101101100: pixel[2:0] = 3'b000;
      14'b00100101101101: pixel[2:0] = 3'b000;
      14'b00100101101110: pixel[2:0] = 3'b000;
      14'b00100101101111: pixel[2:0] = 3'b000;
      14'b00100101110000: pixel[2:0] = 3'b111;
      14'b00100101110001: pixel[2:0] = 3'b111;
      14'b00100101110010: pixel[2:0] = 3'b111;
      14'b00100101110011: pixel[2:0] = 3'b111;
      14'b00100101110100: pixel[2:0] = 3'b111;
      14'b00100101110101: pixel[2:0] = 3'b000;
      14'b00100101110110: pixel[2:0] = 3'b000;
      14'b00100101110111: pixel[2:0] = 3'b000;
      14'b00100101111000: pixel[2:0] = 3'b000;
      14'b00100101111001: pixel[2:0] = 3'b000;
      14'b00100101111010: pixel[2:0] = 3'b000;
      14'b00100101111011: pixel[2:0] = 3'b000;
      14'b00100101111100: pixel[2:0] = 3'b000;
      14'b00100101111101: pixel[2:0] = 3'b111;
      14'b00100101111110: pixel[2:0] = 3'b111;
      14'b00100101111111: pixel[2:0] = 3'b111;
      14'b00100110000000: pixel[2:0] = 3'b111;
      14'b00100110000001: pixel[2:0] = 3'b111;
      14'b00100110000010: pixel[2:0] = 3'b111;
      14'b00100110000011: pixel[2:0] = 3'b000;
      14'b00100110000100: pixel[2:0] = 3'b000;
      14'b00100110000101: pixel[2:0] = 3'b000;
      14'b00100110000110: pixel[2:0] = 3'b000;
      14'b00100110000111: pixel[2:0] = 3'b000;
      14'b00101000000000: pixel[2:0] = 3'b000;
      14'b00101000000001: pixel[2:0] = 3'b000;
      14'b00101000000010: pixel[2:0] = 3'b111;
      14'b00101000000011: pixel[2:0] = 3'b111;
      14'b00101000000100: pixel[2:0] = 3'b111;
      14'b00101000000101: pixel[2:0] = 3'b111;
      14'b00101000000110: pixel[2:0] = 3'b111;
      14'b00101000000111: pixel[2:0] = 3'b000;
      14'b00101000001000: pixel[2:0] = 3'b000;
      14'b00101000001001: pixel[2:0] = 3'b000;
      14'b00101000001010: pixel[2:0] = 3'b000;
      14'b00101000001011: pixel[2:0] = 3'b000;
      14'b00101000001100: pixel[2:0] = 3'b000;
      14'b00101000001101: pixel[2:0] = 3'b000;
      14'b00101000001110: pixel[2:0] = 3'b000;
      14'b00101000001111: pixel[2:0] = 3'b000;
      14'b00101000010000: pixel[2:0] = 3'b111;
      14'b00101000010001: pixel[2:0] = 3'b111;
      14'b00101000010010: pixel[2:0] = 3'b111;
      14'b00101000010011: pixel[2:0] = 3'b111;
      14'b00101000010100: pixel[2:0] = 3'b000;
      14'b00101000010101: pixel[2:0] = 3'b000;
      14'b00101000010110: pixel[2:0] = 3'b000;
      14'b00101000010111: pixel[2:0] = 3'b000;
      14'b00101000011000: pixel[2:0] = 3'b000;
      14'b00101000011001: pixel[2:0] = 3'b111;
      14'b00101000011010: pixel[2:0] = 3'b111;
      14'b00101000011011: pixel[2:0] = 3'b111;
      14'b00101000011100: pixel[2:0] = 3'b111;
      14'b00101000011101: pixel[2:0] = 3'b111;
      14'b00101000011110: pixel[2:0] = 3'b000;
      14'b00101000011111: pixel[2:0] = 3'b000;
      14'b00101000100000: pixel[2:0] = 3'b000;
      14'b00101000100001: pixel[2:0] = 3'b000;
      14'b00101000100010: pixel[2:0] = 3'b000;
      14'b00101000100011: pixel[2:0] = 3'b000;
      14'b00101000100100: pixel[2:0] = 3'b000;
      14'b00101000100101: pixel[2:0] = 3'b000;
      14'b00101000100110: pixel[2:0] = 3'b000;
      14'b00101000100111: pixel[2:0] = 3'b000;
      14'b00101000101000: pixel[2:0] = 3'b000;
      14'b00101000101001: pixel[2:0] = 3'b000;
      14'b00101000101010: pixel[2:0] = 3'b000;
      14'b00101000101011: pixel[2:0] = 3'b000;
      14'b00101000101100: pixel[2:0] = 3'b000;
      14'b00101000101101: pixel[2:0] = 3'b000;
      14'b00101000101110: pixel[2:0] = 3'b000;
      14'b00101000101111: pixel[2:0] = 3'b000;
      14'b00101000110000: pixel[2:0] = 3'b000;
      14'b00101000110001: pixel[2:0] = 3'b000;
      14'b00101000110010: pixel[2:0] = 3'b000;
      14'b00101000110011: pixel[2:0] = 3'b000;
      14'b00101000110100: pixel[2:0] = 3'b111;
      14'b00101000110101: pixel[2:0] = 3'b111;
      14'b00101000110110: pixel[2:0] = 3'b111;
      14'b00101000110111: pixel[2:0] = 3'b111;
      14'b00101000111000: pixel[2:0] = 3'b111;
      14'b00101000111001: pixel[2:0] = 3'b111;
      14'b00101000111010: pixel[2:0] = 3'b111;
      14'b00101000111011: pixel[2:0] = 3'b111;
      14'b00101000111100: pixel[2:0] = 3'b000;
      14'b00101000111101: pixel[2:0] = 3'b000;
      14'b00101000111110: pixel[2:0] = 3'b000;
      14'b00101000111111: pixel[2:0] = 3'b000;
      14'b00101001000000: pixel[2:0] = 3'b000;
      14'b00101001000001: pixel[2:0] = 3'b000;
      14'b00101001000010: pixel[2:0] = 3'b000;
      14'b00101001000011: pixel[2:0] = 3'b000;
      14'b00101001000100: pixel[2:0] = 3'b111;
      14'b00101001000101: pixel[2:0] = 3'b111;
      14'b00101001000110: pixel[2:0] = 3'b111;
      14'b00101001000111: pixel[2:0] = 3'b111;
      14'b00101001001000: pixel[2:0] = 3'b000;
      14'b00101001001001: pixel[2:0] = 3'b000;
      14'b00101001001010: pixel[2:0] = 3'b000;
      14'b00101001001011: pixel[2:0] = 3'b000;
      14'b00101001001100: pixel[2:0] = 3'b000;
      14'b00101001001101: pixel[2:0] = 3'b000;
      14'b00101001001110: pixel[2:0] = 3'b111;
      14'b00101001001111: pixel[2:0] = 3'b111;
      14'b00101001010000: pixel[2:0] = 3'b111;
      14'b00101001010001: pixel[2:0] = 3'b111;
      14'b00101001010010: pixel[2:0] = 3'b111;
      14'b00101001010011: pixel[2:0] = 3'b000;
      14'b00101001010100: pixel[2:0] = 3'b000;
      14'b00101001010101: pixel[2:0] = 3'b000;
      14'b00101001010110: pixel[2:0] = 3'b000;
      14'b00101001010111: pixel[2:0] = 3'b000;
      14'b00101001011000: pixel[2:0] = 3'b000;
      14'b00101001011001: pixel[2:0] = 3'b000;
      14'b00101001011010: pixel[2:0] = 3'b111;
      14'b00101001011011: pixel[2:0] = 3'b111;
      14'b00101001011100: pixel[2:0] = 3'b111;
      14'b00101001011101: pixel[2:0] = 3'b111;
      14'b00101001011110: pixel[2:0] = 3'b111;
      14'b00101001011111: pixel[2:0] = 3'b000;
      14'b00101001100000: pixel[2:0] = 3'b000;
      14'b00101001100001: pixel[2:0] = 3'b000;
      14'b00101001100010: pixel[2:0] = 3'b000;
      14'b00101001100011: pixel[2:0] = 3'b000;
      14'b00101001100100: pixel[2:0] = 3'b000;
      14'b00101001100101: pixel[2:0] = 3'b000;
      14'b00101001100110: pixel[2:0] = 3'b000;
      14'b00101001100111: pixel[2:0] = 3'b000;
      14'b00101001101000: pixel[2:0] = 3'b000;
      14'b00101001101001: pixel[2:0] = 3'b000;
      14'b00101001101010: pixel[2:0] = 3'b000;
      14'b00101001101011: pixel[2:0] = 3'b000;
      14'b00101001101100: pixel[2:0] = 3'b000;
      14'b00101001101101: pixel[2:0] = 3'b000;
      14'b00101001101110: pixel[2:0] = 3'b000;
      14'b00101001101111: pixel[2:0] = 3'b000;
      14'b00101001110000: pixel[2:0] = 3'b111;
      14'b00101001110001: pixel[2:0] = 3'b111;
      14'b00101001110010: pixel[2:0] = 3'b111;
      14'b00101001110011: pixel[2:0] = 3'b111;
      14'b00101001110100: pixel[2:0] = 3'b111;
      14'b00101001110101: pixel[2:0] = 3'b000;
      14'b00101001110110: pixel[2:0] = 3'b000;
      14'b00101001110111: pixel[2:0] = 3'b000;
      14'b00101001111000: pixel[2:0] = 3'b000;
      14'b00101001111001: pixel[2:0] = 3'b000;
      14'b00101001111010: pixel[2:0] = 3'b000;
      14'b00101001111011: pixel[2:0] = 3'b000;
      14'b00101001111100: pixel[2:0] = 3'b000;
      14'b00101001111101: pixel[2:0] = 3'b000;
      14'b00101001111110: pixel[2:0] = 3'b111;
      14'b00101001111111: pixel[2:0] = 3'b111;
      14'b00101010000000: pixel[2:0] = 3'b111;
      14'b00101010000001: pixel[2:0] = 3'b111;
      14'b00101010000010: pixel[2:0] = 3'b111;
      14'b00101010000011: pixel[2:0] = 3'b000;
      14'b00101010000100: pixel[2:0] = 3'b000;
      14'b00101010000101: pixel[2:0] = 3'b000;
      14'b00101010000110: pixel[2:0] = 3'b000;
      14'b00101010000111: pixel[2:0] = 3'b000;
      14'b00101100000000: pixel[2:0] = 3'b000;
      14'b00101100000001: pixel[2:0] = 3'b000;
      14'b00101100000010: pixel[2:0] = 3'b111;
      14'b00101100000011: pixel[2:0] = 3'b111;
      14'b00101100000100: pixel[2:0] = 3'b111;
      14'b00101100000101: pixel[2:0] = 3'b111;
      14'b00101100000110: pixel[2:0] = 3'b111;
      14'b00101100000111: pixel[2:0] = 3'b000;
      14'b00101100001000: pixel[2:0] = 3'b000;
      14'b00101100001001: pixel[2:0] = 3'b000;
      14'b00101100001010: pixel[2:0] = 3'b000;
      14'b00101100001011: pixel[2:0] = 3'b000;
      14'b00101100001100: pixel[2:0] = 3'b000;
      14'b00101100001101: pixel[2:0] = 3'b000;
      14'b00101100001110: pixel[2:0] = 3'b000;
      14'b00101100001111: pixel[2:0] = 3'b000;
      14'b00101100010000: pixel[2:0] = 3'b111;
      14'b00101100010001: pixel[2:0] = 3'b111;
      14'b00101100010010: pixel[2:0] = 3'b111;
      14'b00101100010011: pixel[2:0] = 3'b111;
      14'b00101100010100: pixel[2:0] = 3'b000;
      14'b00101100010101: pixel[2:0] = 3'b000;
      14'b00101100010110: pixel[2:0] = 3'b000;
      14'b00101100010111: pixel[2:0] = 3'b000;
      14'b00101100011000: pixel[2:0] = 3'b000;
      14'b00101100011001: pixel[2:0] = 3'b111;
      14'b00101100011010: pixel[2:0] = 3'b111;
      14'b00101100011011: pixel[2:0] = 3'b111;
      14'b00101100011100: pixel[2:0] = 3'b111;
      14'b00101100011101: pixel[2:0] = 3'b111;
      14'b00101100011110: pixel[2:0] = 3'b000;
      14'b00101100011111: pixel[2:0] = 3'b000;
      14'b00101100100000: pixel[2:0] = 3'b000;
      14'b00101100100001: pixel[2:0] = 3'b000;
      14'b00101100100010: pixel[2:0] = 3'b000;
      14'b00101100100011: pixel[2:0] = 3'b000;
      14'b00101100100100: pixel[2:0] = 3'b000;
      14'b00101100100101: pixel[2:0] = 3'b000;
      14'b00101100100110: pixel[2:0] = 3'b000;
      14'b00101100100111: pixel[2:0] = 3'b000;
      14'b00101100101000: pixel[2:0] = 3'b000;
      14'b00101100101001: pixel[2:0] = 3'b000;
      14'b00101100101010: pixel[2:0] = 3'b000;
      14'b00101100101011: pixel[2:0] = 3'b000;
      14'b00101100101100: pixel[2:0] = 3'b000;
      14'b00101100101101: pixel[2:0] = 3'b000;
      14'b00101100101110: pixel[2:0] = 3'b000;
      14'b00101100101111: pixel[2:0] = 3'b000;
      14'b00101100110000: pixel[2:0] = 3'b000;
      14'b00101100110001: pixel[2:0] = 3'b000;
      14'b00101100110010: pixel[2:0] = 3'b000;
      14'b00101100110011: pixel[2:0] = 3'b000;
      14'b00101100110100: pixel[2:0] = 3'b111;
      14'b00101100110101: pixel[2:0] = 3'b111;
      14'b00101100110110: pixel[2:0] = 3'b111;
      14'b00101100110111: pixel[2:0] = 3'b111;
      14'b00101100111000: pixel[2:0] = 3'b111;
      14'b00101100111001: pixel[2:0] = 3'b111;
      14'b00101100111010: pixel[2:0] = 3'b111;
      14'b00101100111011: pixel[2:0] = 3'b111;
      14'b00101100111100: pixel[2:0] = 3'b000;
      14'b00101100111101: pixel[2:0] = 3'b000;
      14'b00101100111110: pixel[2:0] = 3'b000;
      14'b00101100111111: pixel[2:0] = 3'b000;
      14'b00101101000000: pixel[2:0] = 3'b000;
      14'b00101101000001: pixel[2:0] = 3'b000;
      14'b00101101000010: pixel[2:0] = 3'b000;
      14'b00101101000011: pixel[2:0] = 3'b000;
      14'b00101101000100: pixel[2:0] = 3'b111;
      14'b00101101000101: pixel[2:0] = 3'b111;
      14'b00101101000110: pixel[2:0] = 3'b111;
      14'b00101101000111: pixel[2:0] = 3'b111;
      14'b00101101001000: pixel[2:0] = 3'b111;
      14'b00101101001001: pixel[2:0] = 3'b000;
      14'b00101101001010: pixel[2:0] = 3'b000;
      14'b00101101001011: pixel[2:0] = 3'b000;
      14'b00101101001100: pixel[2:0] = 3'b000;
      14'b00101101001101: pixel[2:0] = 3'b000;
      14'b00101101001110: pixel[2:0] = 3'b111;
      14'b00101101001111: pixel[2:0] = 3'b111;
      14'b00101101010000: pixel[2:0] = 3'b111;
      14'b00101101010001: pixel[2:0] = 3'b111;
      14'b00101101010010: pixel[2:0] = 3'b111;
      14'b00101101010011: pixel[2:0] = 3'b000;
      14'b00101101010100: pixel[2:0] = 3'b000;
      14'b00101101010101: pixel[2:0] = 3'b000;
      14'b00101101010110: pixel[2:0] = 3'b000;
      14'b00101101010111: pixel[2:0] = 3'b000;
      14'b00101101011000: pixel[2:0] = 3'b000;
      14'b00101101011001: pixel[2:0] = 3'b000;
      14'b00101101011010: pixel[2:0] = 3'b111;
      14'b00101101011011: pixel[2:0] = 3'b111;
      14'b00101101011100: pixel[2:0] = 3'b111;
      14'b00101101011101: pixel[2:0] = 3'b111;
      14'b00101101011110: pixel[2:0] = 3'b111;
      14'b00101101011111: pixel[2:0] = 3'b000;
      14'b00101101100000: pixel[2:0] = 3'b000;
      14'b00101101100001: pixel[2:0] = 3'b000;
      14'b00101101100010: pixel[2:0] = 3'b000;
      14'b00101101100011: pixel[2:0] = 3'b000;
      14'b00101101100100: pixel[2:0] = 3'b000;
      14'b00101101100101: pixel[2:0] = 3'b000;
      14'b00101101100110: pixel[2:0] = 3'b000;
      14'b00101101100111: pixel[2:0] = 3'b000;
      14'b00101101101000: pixel[2:0] = 3'b000;
      14'b00101101101001: pixel[2:0] = 3'b000;
      14'b00101101101010: pixel[2:0] = 3'b000;
      14'b00101101101011: pixel[2:0] = 3'b000;
      14'b00101101101100: pixel[2:0] = 3'b000;
      14'b00101101101101: pixel[2:0] = 3'b000;
      14'b00101101101110: pixel[2:0] = 3'b000;
      14'b00101101101111: pixel[2:0] = 3'b000;
      14'b00101101110000: pixel[2:0] = 3'b111;
      14'b00101101110001: pixel[2:0] = 3'b111;
      14'b00101101110010: pixel[2:0] = 3'b111;
      14'b00101101110011: pixel[2:0] = 3'b111;
      14'b00101101110100: pixel[2:0] = 3'b111;
      14'b00101101110101: pixel[2:0] = 3'b000;
      14'b00101101110110: pixel[2:0] = 3'b000;
      14'b00101101110111: pixel[2:0] = 3'b000;
      14'b00101101111000: pixel[2:0] = 3'b000;
      14'b00101101111001: pixel[2:0] = 3'b000;
      14'b00101101111010: pixel[2:0] = 3'b000;
      14'b00101101111011: pixel[2:0] = 3'b000;
      14'b00101101111100: pixel[2:0] = 3'b000;
      14'b00101101111101: pixel[2:0] = 3'b000;
      14'b00101101111110: pixel[2:0] = 3'b111;
      14'b00101101111111: pixel[2:0] = 3'b111;
      14'b00101110000000: pixel[2:0] = 3'b111;
      14'b00101110000001: pixel[2:0] = 3'b111;
      14'b00101110000010: pixel[2:0] = 3'b111;
      14'b00101110000011: pixel[2:0] = 3'b000;
      14'b00101110000100: pixel[2:0] = 3'b000;
      14'b00101110000101: pixel[2:0] = 3'b000;
      14'b00101110000110: pixel[2:0] = 3'b000;
      14'b00101110000111: pixel[2:0] = 3'b000;
      14'b00110000000000: pixel[2:0] = 3'b000;
      14'b00110000000001: pixel[2:0] = 3'b000;
      14'b00110000000010: pixel[2:0] = 3'b111;
      14'b00110000000011: pixel[2:0] = 3'b111;
      14'b00110000000100: pixel[2:0] = 3'b111;
      14'b00110000000101: pixel[2:0] = 3'b111;
      14'b00110000000110: pixel[2:0] = 3'b111;
      14'b00110000000111: pixel[2:0] = 3'b000;
      14'b00110000001000: pixel[2:0] = 3'b000;
      14'b00110000001001: pixel[2:0] = 3'b000;
      14'b00110000001010: pixel[2:0] = 3'b000;
      14'b00110000001011: pixel[2:0] = 3'b000;
      14'b00110000001100: pixel[2:0] = 3'b000;
      14'b00110000001101: pixel[2:0] = 3'b000;
      14'b00110000001110: pixel[2:0] = 3'b000;
      14'b00110000001111: pixel[2:0] = 3'b000;
      14'b00110000010000: pixel[2:0] = 3'b111;
      14'b00110000010001: pixel[2:0] = 3'b111;
      14'b00110000010010: pixel[2:0] = 3'b111;
      14'b00110000010011: pixel[2:0] = 3'b111;
      14'b00110000010100: pixel[2:0] = 3'b000;
      14'b00110000010101: pixel[2:0] = 3'b000;
      14'b00110000010110: pixel[2:0] = 3'b000;
      14'b00110000010111: pixel[2:0] = 3'b000;
      14'b00110000011000: pixel[2:0] = 3'b000;
      14'b00110000011001: pixel[2:0] = 3'b111;
      14'b00110000011010: pixel[2:0] = 3'b111;
      14'b00110000011011: pixel[2:0] = 3'b111;
      14'b00110000011100: pixel[2:0] = 3'b111;
      14'b00110000011101: pixel[2:0] = 3'b111;
      14'b00110000011110: pixel[2:0] = 3'b000;
      14'b00110000011111: pixel[2:0] = 3'b000;
      14'b00110000100000: pixel[2:0] = 3'b000;
      14'b00110000100001: pixel[2:0] = 3'b000;
      14'b00110000100010: pixel[2:0] = 3'b000;
      14'b00110000100011: pixel[2:0] = 3'b000;
      14'b00110000100100: pixel[2:0] = 3'b000;
      14'b00110000100101: pixel[2:0] = 3'b000;
      14'b00110000100110: pixel[2:0] = 3'b000;
      14'b00110000100111: pixel[2:0] = 3'b000;
      14'b00110000101000: pixel[2:0] = 3'b000;
      14'b00110000101001: pixel[2:0] = 3'b000;
      14'b00110000101010: pixel[2:0] = 3'b000;
      14'b00110000101011: pixel[2:0] = 3'b000;
      14'b00110000101100: pixel[2:0] = 3'b000;
      14'b00110000101101: pixel[2:0] = 3'b000;
      14'b00110000101110: pixel[2:0] = 3'b000;
      14'b00110000101111: pixel[2:0] = 3'b000;
      14'b00110000110000: pixel[2:0] = 3'b000;
      14'b00110000110001: pixel[2:0] = 3'b000;
      14'b00110000110010: pixel[2:0] = 3'b000;
      14'b00110000110011: pixel[2:0] = 3'b111;
      14'b00110000110100: pixel[2:0] = 3'b111;
      14'b00110000110101: pixel[2:0] = 3'b111;
      14'b00110000110110: pixel[2:0] = 3'b111;
      14'b00110000110111: pixel[2:0] = 3'b111;
      14'b00110000111000: pixel[2:0] = 3'b111;
      14'b00110000111001: pixel[2:0] = 3'b111;
      14'b00110000111010: pixel[2:0] = 3'b111;
      14'b00110000111011: pixel[2:0] = 3'b111;
      14'b00110000111100: pixel[2:0] = 3'b000;
      14'b00110000111101: pixel[2:0] = 3'b000;
      14'b00110000111110: pixel[2:0] = 3'b000;
      14'b00110000111111: pixel[2:0] = 3'b000;
      14'b00110001000000: pixel[2:0] = 3'b000;
      14'b00110001000001: pixel[2:0] = 3'b000;
      14'b00110001000010: pixel[2:0] = 3'b000;
      14'b00110001000011: pixel[2:0] = 3'b000;
      14'b00110001000100: pixel[2:0] = 3'b111;
      14'b00110001000101: pixel[2:0] = 3'b111;
      14'b00110001000110: pixel[2:0] = 3'b111;
      14'b00110001000111: pixel[2:0] = 3'b111;
      14'b00110001001000: pixel[2:0] = 3'b111;
      14'b00110001001001: pixel[2:0] = 3'b000;
      14'b00110001001010: pixel[2:0] = 3'b000;
      14'b00110001001011: pixel[2:0] = 3'b000;
      14'b00110001001100: pixel[2:0] = 3'b000;
      14'b00110001001101: pixel[2:0] = 3'b000;
      14'b00110001001110: pixel[2:0] = 3'b111;
      14'b00110001001111: pixel[2:0] = 3'b111;
      14'b00110001010000: pixel[2:0] = 3'b111;
      14'b00110001010001: pixel[2:0] = 3'b111;
      14'b00110001010010: pixel[2:0] = 3'b000;
      14'b00110001010011: pixel[2:0] = 3'b000;
      14'b00110001010100: pixel[2:0] = 3'b000;
      14'b00110001010101: pixel[2:0] = 3'b000;
      14'b00110001010110: pixel[2:0] = 3'b000;
      14'b00110001010111: pixel[2:0] = 3'b000;
      14'b00110001011000: pixel[2:0] = 3'b000;
      14'b00110001011001: pixel[2:0] = 3'b000;
      14'b00110001011010: pixel[2:0] = 3'b111;
      14'b00110001011011: pixel[2:0] = 3'b111;
      14'b00110001011100: pixel[2:0] = 3'b111;
      14'b00110001011101: pixel[2:0] = 3'b111;
      14'b00110001011110: pixel[2:0] = 3'b111;
      14'b00110001011111: pixel[2:0] = 3'b000;
      14'b00110001100000: pixel[2:0] = 3'b000;
      14'b00110001100001: pixel[2:0] = 3'b000;
      14'b00110001100010: pixel[2:0] = 3'b000;
      14'b00110001100011: pixel[2:0] = 3'b000;
      14'b00110001100100: pixel[2:0] = 3'b000;
      14'b00110001100101: pixel[2:0] = 3'b000;
      14'b00110001100110: pixel[2:0] = 3'b000;
      14'b00110001100111: pixel[2:0] = 3'b000;
      14'b00110001101000: pixel[2:0] = 3'b000;
      14'b00110001101001: pixel[2:0] = 3'b000;
      14'b00110001101010: pixel[2:0] = 3'b000;
      14'b00110001101011: pixel[2:0] = 3'b000;
      14'b00110001101100: pixel[2:0] = 3'b000;
      14'b00110001101101: pixel[2:0] = 3'b000;
      14'b00110001101110: pixel[2:0] = 3'b000;
      14'b00110001101111: pixel[2:0] = 3'b000;
      14'b00110001110000: pixel[2:0] = 3'b111;
      14'b00110001110001: pixel[2:0] = 3'b111;
      14'b00110001110010: pixel[2:0] = 3'b111;
      14'b00110001110011: pixel[2:0] = 3'b111;
      14'b00110001110100: pixel[2:0] = 3'b111;
      14'b00110001110101: pixel[2:0] = 3'b000;
      14'b00110001110110: pixel[2:0] = 3'b000;
      14'b00110001110111: pixel[2:0] = 3'b000;
      14'b00110001111000: pixel[2:0] = 3'b000;
      14'b00110001111001: pixel[2:0] = 3'b000;
      14'b00110001111010: pixel[2:0] = 3'b000;
      14'b00110001111011: pixel[2:0] = 3'b000;
      14'b00110001111100: pixel[2:0] = 3'b000;
      14'b00110001111101: pixel[2:0] = 3'b000;
      14'b00110001111110: pixel[2:0] = 3'b111;
      14'b00110001111111: pixel[2:0] = 3'b111;
      14'b00110010000000: pixel[2:0] = 3'b111;
      14'b00110010000001: pixel[2:0] = 3'b111;
      14'b00110010000010: pixel[2:0] = 3'b111;
      14'b00110010000011: pixel[2:0] = 3'b000;
      14'b00110010000100: pixel[2:0] = 3'b000;
      14'b00110010000101: pixel[2:0] = 3'b000;
      14'b00110010000110: pixel[2:0] = 3'b000;
      14'b00110010000111: pixel[2:0] = 3'b000;
      14'b00110100000000: pixel[2:0] = 3'b000;
      14'b00110100000001: pixel[2:0] = 3'b000;
      14'b00110100000010: pixel[2:0] = 3'b111;
      14'b00110100000011: pixel[2:0] = 3'b111;
      14'b00110100000100: pixel[2:0] = 3'b111;
      14'b00110100000101: pixel[2:0] = 3'b111;
      14'b00110100000110: pixel[2:0] = 3'b111;
      14'b00110100000111: pixel[2:0] = 3'b000;
      14'b00110100001000: pixel[2:0] = 3'b000;
      14'b00110100001001: pixel[2:0] = 3'b000;
      14'b00110100001010: pixel[2:0] = 3'b000;
      14'b00110100001011: pixel[2:0] = 3'b000;
      14'b00110100001100: pixel[2:0] = 3'b000;
      14'b00110100001101: pixel[2:0] = 3'b000;
      14'b00110100001110: pixel[2:0] = 3'b000;
      14'b00110100001111: pixel[2:0] = 3'b000;
      14'b00110100010000: pixel[2:0] = 3'b111;
      14'b00110100010001: pixel[2:0] = 3'b111;
      14'b00110100010010: pixel[2:0] = 3'b111;
      14'b00110100010011: pixel[2:0] = 3'b111;
      14'b00110100010100: pixel[2:0] = 3'b111;
      14'b00110100010101: pixel[2:0] = 3'b000;
      14'b00110100010110: pixel[2:0] = 3'b000;
      14'b00110100010111: pixel[2:0] = 3'b000;
      14'b00110100011000: pixel[2:0] = 3'b000;
      14'b00110100011001: pixel[2:0] = 3'b111;
      14'b00110100011010: pixel[2:0] = 3'b111;
      14'b00110100011011: pixel[2:0] = 3'b111;
      14'b00110100011100: pixel[2:0] = 3'b111;
      14'b00110100011101: pixel[2:0] = 3'b111;
      14'b00110100011110: pixel[2:0] = 3'b000;
      14'b00110100011111: pixel[2:0] = 3'b000;
      14'b00110100100000: pixel[2:0] = 3'b000;
      14'b00110100100001: pixel[2:0] = 3'b000;
      14'b00110100100010: pixel[2:0] = 3'b000;
      14'b00110100100011: pixel[2:0] = 3'b000;
      14'b00110100100100: pixel[2:0] = 3'b000;
      14'b00110100100101: pixel[2:0] = 3'b000;
      14'b00110100100110: pixel[2:0] = 3'b000;
      14'b00110100100111: pixel[2:0] = 3'b000;
      14'b00110100101000: pixel[2:0] = 3'b000;
      14'b00110100101001: pixel[2:0] = 3'b000;
      14'b00110100101010: pixel[2:0] = 3'b000;
      14'b00110100101011: pixel[2:0] = 3'b000;
      14'b00110100101100: pixel[2:0] = 3'b000;
      14'b00110100101101: pixel[2:0] = 3'b000;
      14'b00110100101110: pixel[2:0] = 3'b000;
      14'b00110100101111: pixel[2:0] = 3'b000;
      14'b00110100110000: pixel[2:0] = 3'b000;
      14'b00110100110001: pixel[2:0] = 3'b000;
      14'b00110100110010: pixel[2:0] = 3'b000;
      14'b00110100110011: pixel[2:0] = 3'b111;
      14'b00110100110100: pixel[2:0] = 3'b111;
      14'b00110100110101: pixel[2:0] = 3'b111;
      14'b00110100110110: pixel[2:0] = 3'b111;
      14'b00110100110111: pixel[2:0] = 3'b111;
      14'b00110100111000: pixel[2:0] = 3'b111;
      14'b00110100111001: pixel[2:0] = 3'b111;
      14'b00110100111010: pixel[2:0] = 3'b111;
      14'b00110100111011: pixel[2:0] = 3'b111;
      14'b00110100111100: pixel[2:0] = 3'b000;
      14'b00110100111101: pixel[2:0] = 3'b000;
      14'b00110100111110: pixel[2:0] = 3'b000;
      14'b00110100111111: pixel[2:0] = 3'b000;
      14'b00110101000000: pixel[2:0] = 3'b000;
      14'b00110101000001: pixel[2:0] = 3'b000;
      14'b00110101000010: pixel[2:0] = 3'b000;
      14'b00110101000011: pixel[2:0] = 3'b000;
      14'b00110101000100: pixel[2:0] = 3'b000;
      14'b00110101000101: pixel[2:0] = 3'b111;
      14'b00110101000110: pixel[2:0] = 3'b111;
      14'b00110101000111: pixel[2:0] = 3'b111;
      14'b00110101001000: pixel[2:0] = 3'b111;
      14'b00110101001001: pixel[2:0] = 3'b000;
      14'b00110101001010: pixel[2:0] = 3'b000;
      14'b00110101001011: pixel[2:0] = 3'b000;
      14'b00110101001100: pixel[2:0] = 3'b000;
      14'b00110101001101: pixel[2:0] = 3'b111;
      14'b00110101001110: pixel[2:0] = 3'b111;
      14'b00110101001111: pixel[2:0] = 3'b111;
      14'b00110101010000: pixel[2:0] = 3'b111;
      14'b00110101010001: pixel[2:0] = 3'b111;
      14'b00110101010010: pixel[2:0] = 3'b000;
      14'b00110101010011: pixel[2:0] = 3'b000;
      14'b00110101010100: pixel[2:0] = 3'b000;
      14'b00110101010101: pixel[2:0] = 3'b000;
      14'b00110101010110: pixel[2:0] = 3'b000;
      14'b00110101010111: pixel[2:0] = 3'b000;
      14'b00110101011000: pixel[2:0] = 3'b000;
      14'b00110101011001: pixel[2:0] = 3'b000;
      14'b00110101011010: pixel[2:0] = 3'b111;
      14'b00110101011011: pixel[2:0] = 3'b111;
      14'b00110101011100: pixel[2:0] = 3'b111;
      14'b00110101011101: pixel[2:0] = 3'b111;
      14'b00110101011110: pixel[2:0] = 3'b111;
      14'b00110101011111: pixel[2:0] = 3'b000;
      14'b00110101100000: pixel[2:0] = 3'b000;
      14'b00110101100001: pixel[2:0] = 3'b000;
      14'b00110101100010: pixel[2:0] = 3'b000;
      14'b00110101100011: pixel[2:0] = 3'b000;
      14'b00110101100100: pixel[2:0] = 3'b000;
      14'b00110101100101: pixel[2:0] = 3'b000;
      14'b00110101100110: pixel[2:0] = 3'b000;
      14'b00110101100111: pixel[2:0] = 3'b000;
      14'b00110101101000: pixel[2:0] = 3'b000;
      14'b00110101101001: pixel[2:0] = 3'b000;
      14'b00110101101010: pixel[2:0] = 3'b000;
      14'b00110101101011: pixel[2:0] = 3'b000;
      14'b00110101101100: pixel[2:0] = 3'b000;
      14'b00110101101101: pixel[2:0] = 3'b000;
      14'b00110101101110: pixel[2:0] = 3'b000;
      14'b00110101101111: pixel[2:0] = 3'b000;
      14'b00110101110000: pixel[2:0] = 3'b111;
      14'b00110101110001: pixel[2:0] = 3'b111;
      14'b00110101110010: pixel[2:0] = 3'b111;
      14'b00110101110011: pixel[2:0] = 3'b111;
      14'b00110101110100: pixel[2:0] = 3'b111;
      14'b00110101110101: pixel[2:0] = 3'b000;
      14'b00110101110110: pixel[2:0] = 3'b000;
      14'b00110101110111: pixel[2:0] = 3'b000;
      14'b00110101111000: pixel[2:0] = 3'b000;
      14'b00110101111001: pixel[2:0] = 3'b000;
      14'b00110101111010: pixel[2:0] = 3'b000;
      14'b00110101111011: pixel[2:0] = 3'b000;
      14'b00110101111100: pixel[2:0] = 3'b000;
      14'b00110101111101: pixel[2:0] = 3'b000;
      14'b00110101111110: pixel[2:0] = 3'b111;
      14'b00110101111111: pixel[2:0] = 3'b111;
      14'b00110110000000: pixel[2:0] = 3'b111;
      14'b00110110000001: pixel[2:0] = 3'b111;
      14'b00110110000010: pixel[2:0] = 3'b111;
      14'b00110110000011: pixel[2:0] = 3'b000;
      14'b00110110000100: pixel[2:0] = 3'b000;
      14'b00110110000101: pixel[2:0] = 3'b000;
      14'b00110110000110: pixel[2:0] = 3'b000;
      14'b00110110000111: pixel[2:0] = 3'b000;
      14'b00111000000000: pixel[2:0] = 3'b000;
      14'b00111000000001: pixel[2:0] = 3'b000;
      14'b00111000000010: pixel[2:0] = 3'b111;
      14'b00111000000011: pixel[2:0] = 3'b111;
      14'b00111000000100: pixel[2:0] = 3'b111;
      14'b00111000000101: pixel[2:0] = 3'b111;
      14'b00111000000110: pixel[2:0] = 3'b111;
      14'b00111000000111: pixel[2:0] = 3'b000;
      14'b00111000001000: pixel[2:0] = 3'b000;
      14'b00111000001001: pixel[2:0] = 3'b000;
      14'b00111000001010: pixel[2:0] = 3'b000;
      14'b00111000001011: pixel[2:0] = 3'b000;
      14'b00111000001100: pixel[2:0] = 3'b000;
      14'b00111000001101: pixel[2:0] = 3'b000;
      14'b00111000001110: pixel[2:0] = 3'b000;
      14'b00111000001111: pixel[2:0] = 3'b000;
      14'b00111000010000: pixel[2:0] = 3'b111;
      14'b00111000010001: pixel[2:0] = 3'b111;
      14'b00111000010010: pixel[2:0] = 3'b111;
      14'b00111000010011: pixel[2:0] = 3'b111;
      14'b00111000010100: pixel[2:0] = 3'b111;
      14'b00111000010101: pixel[2:0] = 3'b000;
      14'b00111000010110: pixel[2:0] = 3'b000;
      14'b00111000010111: pixel[2:0] = 3'b000;
      14'b00111000011000: pixel[2:0] = 3'b000;
      14'b00111000011001: pixel[2:0] = 3'b111;
      14'b00111000011010: pixel[2:0] = 3'b111;
      14'b00111000011011: pixel[2:0] = 3'b111;
      14'b00111000011100: pixel[2:0] = 3'b111;
      14'b00111000011101: pixel[2:0] = 3'b111;
      14'b00111000011110: pixel[2:0] = 3'b000;
      14'b00111000011111: pixel[2:0] = 3'b000;
      14'b00111000100000: pixel[2:0] = 3'b000;
      14'b00111000100001: pixel[2:0] = 3'b000;
      14'b00111000100010: pixel[2:0] = 3'b000;
      14'b00111000100011: pixel[2:0] = 3'b000;
      14'b00111000100100: pixel[2:0] = 3'b000;
      14'b00111000100101: pixel[2:0] = 3'b000;
      14'b00111000100110: pixel[2:0] = 3'b000;
      14'b00111000100111: pixel[2:0] = 3'b000;
      14'b00111000101000: pixel[2:0] = 3'b000;
      14'b00111000101001: pixel[2:0] = 3'b000;
      14'b00111000101010: pixel[2:0] = 3'b000;
      14'b00111000101011: pixel[2:0] = 3'b000;
      14'b00111000101100: pixel[2:0] = 3'b000;
      14'b00111000101101: pixel[2:0] = 3'b000;
      14'b00111000101110: pixel[2:0] = 3'b000;
      14'b00111000101111: pixel[2:0] = 3'b000;
      14'b00111000110000: pixel[2:0] = 3'b000;
      14'b00111000110001: pixel[2:0] = 3'b000;
      14'b00111000110010: pixel[2:0] = 3'b000;
      14'b00111000110011: pixel[2:0] = 3'b111;
      14'b00111000110100: pixel[2:0] = 3'b111;
      14'b00111000110101: pixel[2:0] = 3'b111;
      14'b00111000110110: pixel[2:0] = 3'b111;
      14'b00111000110111: pixel[2:0] = 3'b000;
      14'b00111000111000: pixel[2:0] = 3'b111;
      14'b00111000111001: pixel[2:0] = 3'b111;
      14'b00111000111010: pixel[2:0] = 3'b111;
      14'b00111000111011: pixel[2:0] = 3'b111;
      14'b00111000111100: pixel[2:0] = 3'b111;
      14'b00111000111101: pixel[2:0] = 3'b000;
      14'b00111000111110: pixel[2:0] = 3'b000;
      14'b00111000111111: pixel[2:0] = 3'b000;
      14'b00111001000000: pixel[2:0] = 3'b000;
      14'b00111001000001: pixel[2:0] = 3'b000;
      14'b00111001000010: pixel[2:0] = 3'b000;
      14'b00111001000011: pixel[2:0] = 3'b000;
      14'b00111001000100: pixel[2:0] = 3'b000;
      14'b00111001000101: pixel[2:0] = 3'b111;
      14'b00111001000110: pixel[2:0] = 3'b111;
      14'b00111001000111: pixel[2:0] = 3'b111;
      14'b00111001001000: pixel[2:0] = 3'b111;
      14'b00111001001001: pixel[2:0] = 3'b111;
      14'b00111001001010: pixel[2:0] = 3'b000;
      14'b00111001001011: pixel[2:0] = 3'b000;
      14'b00111001001100: pixel[2:0] = 3'b000;
      14'b00111001001101: pixel[2:0] = 3'b111;
      14'b00111001001110: pixel[2:0] = 3'b111;
      14'b00111001001111: pixel[2:0] = 3'b111;
      14'b00111001010000: pixel[2:0] = 3'b111;
      14'b00111001010001: pixel[2:0] = 3'b111;
      14'b00111001010010: pixel[2:0] = 3'b000;
      14'b00111001010011: pixel[2:0] = 3'b000;
      14'b00111001010100: pixel[2:0] = 3'b000;
      14'b00111001010101: pixel[2:0] = 3'b000;
      14'b00111001010110: pixel[2:0] = 3'b000;
      14'b00111001010111: pixel[2:0] = 3'b000;
      14'b00111001011000: pixel[2:0] = 3'b000;
      14'b00111001011001: pixel[2:0] = 3'b000;
      14'b00111001011010: pixel[2:0] = 3'b111;
      14'b00111001011011: pixel[2:0] = 3'b111;
      14'b00111001011100: pixel[2:0] = 3'b111;
      14'b00111001011101: pixel[2:0] = 3'b111;
      14'b00111001011110: pixel[2:0] = 3'b111;
      14'b00111001011111: pixel[2:0] = 3'b000;
      14'b00111001100000: pixel[2:0] = 3'b000;
      14'b00111001100001: pixel[2:0] = 3'b000;
      14'b00111001100010: pixel[2:0] = 3'b000;
      14'b00111001100011: pixel[2:0] = 3'b000;
      14'b00111001100100: pixel[2:0] = 3'b000;
      14'b00111001100101: pixel[2:0] = 3'b000;
      14'b00111001100110: pixel[2:0] = 3'b000;
      14'b00111001100111: pixel[2:0] = 3'b000;
      14'b00111001101000: pixel[2:0] = 3'b000;
      14'b00111001101001: pixel[2:0] = 3'b000;
      14'b00111001101010: pixel[2:0] = 3'b000;
      14'b00111001101011: pixel[2:0] = 3'b000;
      14'b00111001101100: pixel[2:0] = 3'b000;
      14'b00111001101101: pixel[2:0] = 3'b000;
      14'b00111001101110: pixel[2:0] = 3'b000;
      14'b00111001101111: pixel[2:0] = 3'b000;
      14'b00111001110000: pixel[2:0] = 3'b111;
      14'b00111001110001: pixel[2:0] = 3'b111;
      14'b00111001110010: pixel[2:0] = 3'b111;
      14'b00111001110011: pixel[2:0] = 3'b111;
      14'b00111001110100: pixel[2:0] = 3'b111;
      14'b00111001110101: pixel[2:0] = 3'b000;
      14'b00111001110110: pixel[2:0] = 3'b000;
      14'b00111001110111: pixel[2:0] = 3'b000;
      14'b00111001111000: pixel[2:0] = 3'b000;
      14'b00111001111001: pixel[2:0] = 3'b000;
      14'b00111001111010: pixel[2:0] = 3'b000;
      14'b00111001111011: pixel[2:0] = 3'b000;
      14'b00111001111100: pixel[2:0] = 3'b000;
      14'b00111001111101: pixel[2:0] = 3'b000;
      14'b00111001111110: pixel[2:0] = 3'b111;
      14'b00111001111111: pixel[2:0] = 3'b111;
      14'b00111010000000: pixel[2:0] = 3'b111;
      14'b00111010000001: pixel[2:0] = 3'b111;
      14'b00111010000010: pixel[2:0] = 3'b111;
      14'b00111010000011: pixel[2:0] = 3'b000;
      14'b00111010000100: pixel[2:0] = 3'b000;
      14'b00111010000101: pixel[2:0] = 3'b000;
      14'b00111010000110: pixel[2:0] = 3'b000;
      14'b00111010000111: pixel[2:0] = 3'b000;
      14'b00111100000000: pixel[2:0] = 3'b000;
      14'b00111100000001: pixel[2:0] = 3'b000;
      14'b00111100000010: pixel[2:0] = 3'b111;
      14'b00111100000011: pixel[2:0] = 3'b111;
      14'b00111100000100: pixel[2:0] = 3'b111;
      14'b00111100000101: pixel[2:0] = 3'b111;
      14'b00111100000110: pixel[2:0] = 3'b111;
      14'b00111100000111: pixel[2:0] = 3'b000;
      14'b00111100001000: pixel[2:0] = 3'b000;
      14'b00111100001001: pixel[2:0] = 3'b000;
      14'b00111100001010: pixel[2:0] = 3'b000;
      14'b00111100001011: pixel[2:0] = 3'b000;
      14'b00111100001100: pixel[2:0] = 3'b000;
      14'b00111100001101: pixel[2:0] = 3'b000;
      14'b00111100001110: pixel[2:0] = 3'b000;
      14'b00111100001111: pixel[2:0] = 3'b000;
      14'b00111100010000: pixel[2:0] = 3'b111;
      14'b00111100010001: pixel[2:0] = 3'b111;
      14'b00111100010010: pixel[2:0] = 3'b111;
      14'b00111100010011: pixel[2:0] = 3'b111;
      14'b00111100010100: pixel[2:0] = 3'b111;
      14'b00111100010101: pixel[2:0] = 3'b000;
      14'b00111100010110: pixel[2:0] = 3'b000;
      14'b00111100010111: pixel[2:0] = 3'b000;
      14'b00111100011000: pixel[2:0] = 3'b000;
      14'b00111100011001: pixel[2:0] = 3'b111;
      14'b00111100011010: pixel[2:0] = 3'b111;
      14'b00111100011011: pixel[2:0] = 3'b111;
      14'b00111100011100: pixel[2:0] = 3'b111;
      14'b00111100011101: pixel[2:0] = 3'b111;
      14'b00111100011110: pixel[2:0] = 3'b000;
      14'b00111100011111: pixel[2:0] = 3'b000;
      14'b00111100100000: pixel[2:0] = 3'b000;
      14'b00111100100001: pixel[2:0] = 3'b000;
      14'b00111100100010: pixel[2:0] = 3'b000;
      14'b00111100100011: pixel[2:0] = 3'b000;
      14'b00111100100100: pixel[2:0] = 3'b000;
      14'b00111100100101: pixel[2:0] = 3'b000;
      14'b00111100100110: pixel[2:0] = 3'b000;
      14'b00111100100111: pixel[2:0] = 3'b000;
      14'b00111100101000: pixel[2:0] = 3'b000;
      14'b00111100101001: pixel[2:0] = 3'b000;
      14'b00111100101010: pixel[2:0] = 3'b000;
      14'b00111100101011: pixel[2:0] = 3'b000;
      14'b00111100101100: pixel[2:0] = 3'b000;
      14'b00111100101101: pixel[2:0] = 3'b000;
      14'b00111100101110: pixel[2:0] = 3'b000;
      14'b00111100101111: pixel[2:0] = 3'b000;
      14'b00111100110000: pixel[2:0] = 3'b000;
      14'b00111100110001: pixel[2:0] = 3'b000;
      14'b00111100110010: pixel[2:0] = 3'b000;
      14'b00111100110011: pixel[2:0] = 3'b111;
      14'b00111100110100: pixel[2:0] = 3'b111;
      14'b00111100110101: pixel[2:0] = 3'b111;
      14'b00111100110110: pixel[2:0] = 3'b111;
      14'b00111100110111: pixel[2:0] = 3'b000;
      14'b00111100111000: pixel[2:0] = 3'b000;
      14'b00111100111001: pixel[2:0] = 3'b111;
      14'b00111100111010: pixel[2:0] = 3'b111;
      14'b00111100111011: pixel[2:0] = 3'b111;
      14'b00111100111100: pixel[2:0] = 3'b111;
      14'b00111100111101: pixel[2:0] = 3'b000;
      14'b00111100111110: pixel[2:0] = 3'b000;
      14'b00111100111111: pixel[2:0] = 3'b000;
      14'b00111101000000: pixel[2:0] = 3'b000;
      14'b00111101000001: pixel[2:0] = 3'b000;
      14'b00111101000010: pixel[2:0] = 3'b000;
      14'b00111101000011: pixel[2:0] = 3'b000;
      14'b00111101000100: pixel[2:0] = 3'b000;
      14'b00111101000101: pixel[2:0] = 3'b111;
      14'b00111101000110: pixel[2:0] = 3'b111;
      14'b00111101000111: pixel[2:0] = 3'b111;
      14'b00111101001000: pixel[2:0] = 3'b111;
      14'b00111101001001: pixel[2:0] = 3'b111;
      14'b00111101001010: pixel[2:0] = 3'b000;
      14'b00111101001011: pixel[2:0] = 3'b000;
      14'b00111101001100: pixel[2:0] = 3'b000;
      14'b00111101001101: pixel[2:0] = 3'b111;
      14'b00111101001110: pixel[2:0] = 3'b111;
      14'b00111101001111: pixel[2:0] = 3'b111;
      14'b00111101010000: pixel[2:0] = 3'b111;
      14'b00111101010001: pixel[2:0] = 3'b000;
      14'b00111101010010: pixel[2:0] = 3'b000;
      14'b00111101010011: pixel[2:0] = 3'b000;
      14'b00111101010100: pixel[2:0] = 3'b000;
      14'b00111101010101: pixel[2:0] = 3'b000;
      14'b00111101010110: pixel[2:0] = 3'b000;
      14'b00111101010111: pixel[2:0] = 3'b000;
      14'b00111101011000: pixel[2:0] = 3'b000;
      14'b00111101011001: pixel[2:0] = 3'b000;
      14'b00111101011010: pixel[2:0] = 3'b111;
      14'b00111101011011: pixel[2:0] = 3'b111;
      14'b00111101011100: pixel[2:0] = 3'b111;
      14'b00111101011101: pixel[2:0] = 3'b111;
      14'b00111101011110: pixel[2:0] = 3'b111;
      14'b00111101011111: pixel[2:0] = 3'b000;
      14'b00111101100000: pixel[2:0] = 3'b000;
      14'b00111101100001: pixel[2:0] = 3'b000;
      14'b00111101100010: pixel[2:0] = 3'b000;
      14'b00111101100011: pixel[2:0] = 3'b000;
      14'b00111101100100: pixel[2:0] = 3'b000;
      14'b00111101100101: pixel[2:0] = 3'b000;
      14'b00111101100110: pixel[2:0] = 3'b000;
      14'b00111101100111: pixel[2:0] = 3'b000;
      14'b00111101101000: pixel[2:0] = 3'b000;
      14'b00111101101001: pixel[2:0] = 3'b000;
      14'b00111101101010: pixel[2:0] = 3'b000;
      14'b00111101101011: pixel[2:0] = 3'b000;
      14'b00111101101100: pixel[2:0] = 3'b000;
      14'b00111101101101: pixel[2:0] = 3'b000;
      14'b00111101101110: pixel[2:0] = 3'b000;
      14'b00111101101111: pixel[2:0] = 3'b000;
      14'b00111101110000: pixel[2:0] = 3'b111;
      14'b00111101110001: pixel[2:0] = 3'b111;
      14'b00111101110010: pixel[2:0] = 3'b111;
      14'b00111101110011: pixel[2:0] = 3'b111;
      14'b00111101110100: pixel[2:0] = 3'b111;
      14'b00111101110101: pixel[2:0] = 3'b000;
      14'b00111101110110: pixel[2:0] = 3'b000;
      14'b00111101110111: pixel[2:0] = 3'b000;
      14'b00111101111000: pixel[2:0] = 3'b000;
      14'b00111101111001: pixel[2:0] = 3'b000;
      14'b00111101111010: pixel[2:0] = 3'b000;
      14'b00111101111011: pixel[2:0] = 3'b000;
      14'b00111101111100: pixel[2:0] = 3'b000;
      14'b00111101111101: pixel[2:0] = 3'b000;
      14'b00111101111110: pixel[2:0] = 3'b111;
      14'b00111101111111: pixel[2:0] = 3'b111;
      14'b00111110000000: pixel[2:0] = 3'b111;
      14'b00111110000001: pixel[2:0] = 3'b111;
      14'b00111110000010: pixel[2:0] = 3'b111;
      14'b00111110000011: pixel[2:0] = 3'b000;
      14'b00111110000100: pixel[2:0] = 3'b000;
      14'b00111110000101: pixel[2:0] = 3'b000;
      14'b00111110000110: pixel[2:0] = 3'b000;
      14'b00111110000111: pixel[2:0] = 3'b000;
      14'b01000000000000: pixel[2:0] = 3'b000;
      14'b01000000000001: pixel[2:0] = 3'b000;
      14'b01000000000010: pixel[2:0] = 3'b111;
      14'b01000000000011: pixel[2:0] = 3'b111;
      14'b01000000000100: pixel[2:0] = 3'b111;
      14'b01000000000101: pixel[2:0] = 3'b111;
      14'b01000000000110: pixel[2:0] = 3'b111;
      14'b01000000000111: pixel[2:0] = 3'b000;
      14'b01000000001000: pixel[2:0] = 3'b000;
      14'b01000000001001: pixel[2:0] = 3'b000;
      14'b01000000001010: pixel[2:0] = 3'b000;
      14'b01000000001011: pixel[2:0] = 3'b000;
      14'b01000000001100: pixel[2:0] = 3'b000;
      14'b01000000001101: pixel[2:0] = 3'b000;
      14'b01000000001110: pixel[2:0] = 3'b000;
      14'b01000000001111: pixel[2:0] = 3'b000;
      14'b01000000010000: pixel[2:0] = 3'b111;
      14'b01000000010001: pixel[2:0] = 3'b111;
      14'b01000000010010: pixel[2:0] = 3'b111;
      14'b01000000010011: pixel[2:0] = 3'b111;
      14'b01000000010100: pixel[2:0] = 3'b000;
      14'b01000000010101: pixel[2:0] = 3'b000;
      14'b01000000010110: pixel[2:0] = 3'b000;
      14'b01000000010111: pixel[2:0] = 3'b000;
      14'b01000000011000: pixel[2:0] = 3'b000;
      14'b01000000011001: pixel[2:0] = 3'b111;
      14'b01000000011010: pixel[2:0] = 3'b111;
      14'b01000000011011: pixel[2:0] = 3'b111;
      14'b01000000011100: pixel[2:0] = 3'b111;
      14'b01000000011101: pixel[2:0] = 3'b111;
      14'b01000000011110: pixel[2:0] = 3'b000;
      14'b01000000011111: pixel[2:0] = 3'b000;
      14'b01000000100000: pixel[2:0] = 3'b000;
      14'b01000000100001: pixel[2:0] = 3'b000;
      14'b01000000100010: pixel[2:0] = 3'b000;
      14'b01000000100011: pixel[2:0] = 3'b000;
      14'b01000000100100: pixel[2:0] = 3'b000;
      14'b01000000100101: pixel[2:0] = 3'b000;
      14'b01000000100110: pixel[2:0] = 3'b000;
      14'b01000000100111: pixel[2:0] = 3'b000;
      14'b01000000101000: pixel[2:0] = 3'b000;
      14'b01000000101001: pixel[2:0] = 3'b000;
      14'b01000000101010: pixel[2:0] = 3'b000;
      14'b01000000101011: pixel[2:0] = 3'b000;
      14'b01000000101100: pixel[2:0] = 3'b000;
      14'b01000000101101: pixel[2:0] = 3'b000;
      14'b01000000101110: pixel[2:0] = 3'b000;
      14'b01000000101111: pixel[2:0] = 3'b000;
      14'b01000000110000: pixel[2:0] = 3'b000;
      14'b01000000110001: pixel[2:0] = 3'b000;
      14'b01000000110010: pixel[2:0] = 3'b000;
      14'b01000000110011: pixel[2:0] = 3'b111;
      14'b01000000110100: pixel[2:0] = 3'b111;
      14'b01000000110101: pixel[2:0] = 3'b111;
      14'b01000000110110: pixel[2:0] = 3'b111;
      14'b01000000110111: pixel[2:0] = 3'b000;
      14'b01000000111000: pixel[2:0] = 3'b000;
      14'b01000000111001: pixel[2:0] = 3'b111;
      14'b01000000111010: pixel[2:0] = 3'b111;
      14'b01000000111011: pixel[2:0] = 3'b111;
      14'b01000000111100: pixel[2:0] = 3'b111;
      14'b01000000111101: pixel[2:0] = 3'b000;
      14'b01000000111110: pixel[2:0] = 3'b000;
      14'b01000000111111: pixel[2:0] = 3'b000;
      14'b01000001000000: pixel[2:0] = 3'b000;
      14'b01000001000001: pixel[2:0] = 3'b000;
      14'b01000001000010: pixel[2:0] = 3'b000;
      14'b01000001000011: pixel[2:0] = 3'b000;
      14'b01000001000100: pixel[2:0] = 3'b000;
      14'b01000001000101: pixel[2:0] = 3'b000;
      14'b01000001000110: pixel[2:0] = 3'b111;
      14'b01000001000111: pixel[2:0] = 3'b111;
      14'b01000001001000: pixel[2:0] = 3'b111;
      14'b01000001001001: pixel[2:0] = 3'b111;
      14'b01000001001010: pixel[2:0] = 3'b000;
      14'b01000001001011: pixel[2:0] = 3'b000;
      14'b01000001001100: pixel[2:0] = 3'b111;
      14'b01000001001101: pixel[2:0] = 3'b111;
      14'b01000001001110: pixel[2:0] = 3'b111;
      14'b01000001001111: pixel[2:0] = 3'b111;
      14'b01000001010000: pixel[2:0] = 3'b111;
      14'b01000001010001: pixel[2:0] = 3'b000;
      14'b01000001010010: pixel[2:0] = 3'b000;
      14'b01000001010011: pixel[2:0] = 3'b000;
      14'b01000001010100: pixel[2:0] = 3'b000;
      14'b01000001010101: pixel[2:0] = 3'b000;
      14'b01000001010110: pixel[2:0] = 3'b000;
      14'b01000001010111: pixel[2:0] = 3'b000;
      14'b01000001011000: pixel[2:0] = 3'b000;
      14'b01000001011001: pixel[2:0] = 3'b000;
      14'b01000001011010: pixel[2:0] = 3'b111;
      14'b01000001011011: pixel[2:0] = 3'b111;
      14'b01000001011100: pixel[2:0] = 3'b111;
      14'b01000001011101: pixel[2:0] = 3'b111;
      14'b01000001011110: pixel[2:0] = 3'b111;
      14'b01000001011111: pixel[2:0] = 3'b000;
      14'b01000001100000: pixel[2:0] = 3'b000;
      14'b01000001100001: pixel[2:0] = 3'b000;
      14'b01000001100010: pixel[2:0] = 3'b000;
      14'b01000001100011: pixel[2:0] = 3'b000;
      14'b01000001100100: pixel[2:0] = 3'b000;
      14'b01000001100101: pixel[2:0] = 3'b000;
      14'b01000001100110: pixel[2:0] = 3'b000;
      14'b01000001100111: pixel[2:0] = 3'b000;
      14'b01000001101000: pixel[2:0] = 3'b000;
      14'b01000001101001: pixel[2:0] = 3'b000;
      14'b01000001101010: pixel[2:0] = 3'b000;
      14'b01000001101011: pixel[2:0] = 3'b000;
      14'b01000001101100: pixel[2:0] = 3'b000;
      14'b01000001101101: pixel[2:0] = 3'b000;
      14'b01000001101110: pixel[2:0] = 3'b000;
      14'b01000001101111: pixel[2:0] = 3'b000;
      14'b01000001110000: pixel[2:0] = 3'b111;
      14'b01000001110001: pixel[2:0] = 3'b111;
      14'b01000001110010: pixel[2:0] = 3'b111;
      14'b01000001110011: pixel[2:0] = 3'b111;
      14'b01000001110100: pixel[2:0] = 3'b111;
      14'b01000001110101: pixel[2:0] = 3'b000;
      14'b01000001110110: pixel[2:0] = 3'b000;
      14'b01000001110111: pixel[2:0] = 3'b000;
      14'b01000001111000: pixel[2:0] = 3'b000;
      14'b01000001111001: pixel[2:0] = 3'b000;
      14'b01000001111010: pixel[2:0] = 3'b000;
      14'b01000001111011: pixel[2:0] = 3'b000;
      14'b01000001111100: pixel[2:0] = 3'b000;
      14'b01000001111101: pixel[2:0] = 3'b000;
      14'b01000001111110: pixel[2:0] = 3'b111;
      14'b01000001111111: pixel[2:0] = 3'b111;
      14'b01000010000000: pixel[2:0] = 3'b111;
      14'b01000010000001: pixel[2:0] = 3'b111;
      14'b01000010000010: pixel[2:0] = 3'b111;
      14'b01000010000011: pixel[2:0] = 3'b000;
      14'b01000010000100: pixel[2:0] = 3'b000;
      14'b01000010000101: pixel[2:0] = 3'b000;
      14'b01000010000110: pixel[2:0] = 3'b000;
      14'b01000010000111: pixel[2:0] = 3'b000;
      14'b01000100000000: pixel[2:0] = 3'b000;
      14'b01000100000001: pixel[2:0] = 3'b000;
      14'b01000100000010: pixel[2:0] = 3'b111;
      14'b01000100000011: pixel[2:0] = 3'b111;
      14'b01000100000100: pixel[2:0] = 3'b111;
      14'b01000100000101: pixel[2:0] = 3'b111;
      14'b01000100000110: pixel[2:0] = 3'b111;
      14'b01000100000111: pixel[2:0] = 3'b000;
      14'b01000100001000: pixel[2:0] = 3'b000;
      14'b01000100001001: pixel[2:0] = 3'b000;
      14'b01000100001010: pixel[2:0] = 3'b000;
      14'b01000100001011: pixel[2:0] = 3'b000;
      14'b01000100001100: pixel[2:0] = 3'b000;
      14'b01000100001101: pixel[2:0] = 3'b000;
      14'b01000100001110: pixel[2:0] = 3'b000;
      14'b01000100001111: pixel[2:0] = 3'b000;
      14'b01000100010000: pixel[2:0] = 3'b111;
      14'b01000100010001: pixel[2:0] = 3'b111;
      14'b01000100010010: pixel[2:0] = 3'b111;
      14'b01000100010011: pixel[2:0] = 3'b111;
      14'b01000100010100: pixel[2:0] = 3'b000;
      14'b01000100010101: pixel[2:0] = 3'b000;
      14'b01000100010110: pixel[2:0] = 3'b000;
      14'b01000100010111: pixel[2:0] = 3'b000;
      14'b01000100011000: pixel[2:0] = 3'b000;
      14'b01000100011001: pixel[2:0] = 3'b111;
      14'b01000100011010: pixel[2:0] = 3'b111;
      14'b01000100011011: pixel[2:0] = 3'b111;
      14'b01000100011100: pixel[2:0] = 3'b111;
      14'b01000100011101: pixel[2:0] = 3'b111;
      14'b01000100011110: pixel[2:0] = 3'b000;
      14'b01000100011111: pixel[2:0] = 3'b000;
      14'b01000100100000: pixel[2:0] = 3'b000;
      14'b01000100100001: pixel[2:0] = 3'b000;
      14'b01000100100010: pixel[2:0] = 3'b000;
      14'b01000100100011: pixel[2:0] = 3'b000;
      14'b01000100100100: pixel[2:0] = 3'b000;
      14'b01000100100101: pixel[2:0] = 3'b000;
      14'b01000100100110: pixel[2:0] = 3'b000;
      14'b01000100100111: pixel[2:0] = 3'b000;
      14'b01000100101000: pixel[2:0] = 3'b000;
      14'b01000100101001: pixel[2:0] = 3'b000;
      14'b01000100101010: pixel[2:0] = 3'b000;
      14'b01000100101011: pixel[2:0] = 3'b000;
      14'b01000100101100: pixel[2:0] = 3'b000;
      14'b01000100101101: pixel[2:0] = 3'b000;
      14'b01000100101110: pixel[2:0] = 3'b000;
      14'b01000100101111: pixel[2:0] = 3'b000;
      14'b01000100110000: pixel[2:0] = 3'b000;
      14'b01000100110001: pixel[2:0] = 3'b000;
      14'b01000100110010: pixel[2:0] = 3'b111;
      14'b01000100110011: pixel[2:0] = 3'b111;
      14'b01000100110100: pixel[2:0] = 3'b111;
      14'b01000100110101: pixel[2:0] = 3'b111;
      14'b01000100110110: pixel[2:0] = 3'b000;
      14'b01000100110111: pixel[2:0] = 3'b000;
      14'b01000100111000: pixel[2:0] = 3'b000;
      14'b01000100111001: pixel[2:0] = 3'b111;
      14'b01000100111010: pixel[2:0] = 3'b111;
      14'b01000100111011: pixel[2:0] = 3'b111;
      14'b01000100111100: pixel[2:0] = 3'b111;
      14'b01000100111101: pixel[2:0] = 3'b000;
      14'b01000100111110: pixel[2:0] = 3'b000;
      14'b01000100111111: pixel[2:0] = 3'b000;
      14'b01000101000000: pixel[2:0] = 3'b000;
      14'b01000101000001: pixel[2:0] = 3'b000;
      14'b01000101000010: pixel[2:0] = 3'b000;
      14'b01000101000011: pixel[2:0] = 3'b000;
      14'b01000101000100: pixel[2:0] = 3'b000;
      14'b01000101000101: pixel[2:0] = 3'b000;
      14'b01000101000110: pixel[2:0] = 3'b111;
      14'b01000101000111: pixel[2:0] = 3'b111;
      14'b01000101001000: pixel[2:0] = 3'b111;
      14'b01000101001001: pixel[2:0] = 3'b111;
      14'b01000101001010: pixel[2:0] = 3'b000;
      14'b01000101001011: pixel[2:0] = 3'b000;
      14'b01000101001100: pixel[2:0] = 3'b111;
      14'b01000101001101: pixel[2:0] = 3'b111;
      14'b01000101001110: pixel[2:0] = 3'b111;
      14'b01000101001111: pixel[2:0] = 3'b111;
      14'b01000101010000: pixel[2:0] = 3'b000;
      14'b01000101010001: pixel[2:0] = 3'b000;
      14'b01000101010010: pixel[2:0] = 3'b000;
      14'b01000101010011: pixel[2:0] = 3'b000;
      14'b01000101010100: pixel[2:0] = 3'b000;
      14'b01000101010101: pixel[2:0] = 3'b000;
      14'b01000101010110: pixel[2:0] = 3'b000;
      14'b01000101010111: pixel[2:0] = 3'b000;
      14'b01000101011000: pixel[2:0] = 3'b000;
      14'b01000101011001: pixel[2:0] = 3'b000;
      14'b01000101011010: pixel[2:0] = 3'b111;
      14'b01000101011011: pixel[2:0] = 3'b111;
      14'b01000101011100: pixel[2:0] = 3'b111;
      14'b01000101011101: pixel[2:0] = 3'b111;
      14'b01000101011110: pixel[2:0] = 3'b111;
      14'b01000101011111: pixel[2:0] = 3'b000;
      14'b01000101100000: pixel[2:0] = 3'b000;
      14'b01000101100001: pixel[2:0] = 3'b000;
      14'b01000101100010: pixel[2:0] = 3'b000;
      14'b01000101100011: pixel[2:0] = 3'b000;
      14'b01000101100100: pixel[2:0] = 3'b000;
      14'b01000101100101: pixel[2:0] = 3'b000;
      14'b01000101100110: pixel[2:0] = 3'b000;
      14'b01000101100111: pixel[2:0] = 3'b000;
      14'b01000101101000: pixel[2:0] = 3'b000;
      14'b01000101101001: pixel[2:0] = 3'b000;
      14'b01000101101010: pixel[2:0] = 3'b000;
      14'b01000101101011: pixel[2:0] = 3'b000;
      14'b01000101101100: pixel[2:0] = 3'b000;
      14'b01000101101101: pixel[2:0] = 3'b000;
      14'b01000101101110: pixel[2:0] = 3'b000;
      14'b01000101101111: pixel[2:0] = 3'b000;
      14'b01000101110000: pixel[2:0] = 3'b111;
      14'b01000101110001: pixel[2:0] = 3'b111;
      14'b01000101110010: pixel[2:0] = 3'b111;
      14'b01000101110011: pixel[2:0] = 3'b111;
      14'b01000101110100: pixel[2:0] = 3'b111;
      14'b01000101110101: pixel[2:0] = 3'b000;
      14'b01000101110110: pixel[2:0] = 3'b000;
      14'b01000101110111: pixel[2:0] = 3'b000;
      14'b01000101111000: pixel[2:0] = 3'b000;
      14'b01000101111001: pixel[2:0] = 3'b000;
      14'b01000101111010: pixel[2:0] = 3'b000;
      14'b01000101111011: pixel[2:0] = 3'b000;
      14'b01000101111100: pixel[2:0] = 3'b000;
      14'b01000101111101: pixel[2:0] = 3'b000;
      14'b01000101111110: pixel[2:0] = 3'b111;
      14'b01000101111111: pixel[2:0] = 3'b111;
      14'b01000110000000: pixel[2:0] = 3'b111;
      14'b01000110000001: pixel[2:0] = 3'b111;
      14'b01000110000010: pixel[2:0] = 3'b111;
      14'b01000110000011: pixel[2:0] = 3'b000;
      14'b01000110000100: pixel[2:0] = 3'b000;
      14'b01000110000101: pixel[2:0] = 3'b000;
      14'b01000110000110: pixel[2:0] = 3'b000;
      14'b01000110000111: pixel[2:0] = 3'b000;
      14'b01001000000000: pixel[2:0] = 3'b000;
      14'b01001000000001: pixel[2:0] = 3'b000;
      14'b01001000000010: pixel[2:0] = 3'b111;
      14'b01001000000011: pixel[2:0] = 3'b111;
      14'b01001000000100: pixel[2:0] = 3'b111;
      14'b01001000000101: pixel[2:0] = 3'b111;
      14'b01001000000110: pixel[2:0] = 3'b111;
      14'b01001000000111: pixel[2:0] = 3'b000;
      14'b01001000001000: pixel[2:0] = 3'b000;
      14'b01001000001001: pixel[2:0] = 3'b000;
      14'b01001000001010: pixel[2:0] = 3'b000;
      14'b01001000001011: pixel[2:0] = 3'b000;
      14'b01001000001100: pixel[2:0] = 3'b000;
      14'b01001000001101: pixel[2:0] = 3'b000;
      14'b01001000001110: pixel[2:0] = 3'b000;
      14'b01001000001111: pixel[2:0] = 3'b000;
      14'b01001000010000: pixel[2:0] = 3'b111;
      14'b01001000010001: pixel[2:0] = 3'b111;
      14'b01001000010010: pixel[2:0] = 3'b111;
      14'b01001000010011: pixel[2:0] = 3'b111;
      14'b01001000010100: pixel[2:0] = 3'b000;
      14'b01001000010101: pixel[2:0] = 3'b000;
      14'b01001000010110: pixel[2:0] = 3'b000;
      14'b01001000010111: pixel[2:0] = 3'b000;
      14'b01001000011000: pixel[2:0] = 3'b000;
      14'b01001000011001: pixel[2:0] = 3'b111;
      14'b01001000011010: pixel[2:0] = 3'b111;
      14'b01001000011011: pixel[2:0] = 3'b111;
      14'b01001000011100: pixel[2:0] = 3'b111;
      14'b01001000011101: pixel[2:0] = 3'b111;
      14'b01001000011110: pixel[2:0] = 3'b000;
      14'b01001000011111: pixel[2:0] = 3'b000;
      14'b01001000100000: pixel[2:0] = 3'b000;
      14'b01001000100001: pixel[2:0] = 3'b000;
      14'b01001000100010: pixel[2:0] = 3'b000;
      14'b01001000100011: pixel[2:0] = 3'b000;
      14'b01001000100100: pixel[2:0] = 3'b000;
      14'b01001000100101: pixel[2:0] = 3'b000;
      14'b01001000100110: pixel[2:0] = 3'b000;
      14'b01001000100111: pixel[2:0] = 3'b000;
      14'b01001000101000: pixel[2:0] = 3'b000;
      14'b01001000101001: pixel[2:0] = 3'b000;
      14'b01001000101010: pixel[2:0] = 3'b000;
      14'b01001000101011: pixel[2:0] = 3'b000;
      14'b01001000101100: pixel[2:0] = 3'b000;
      14'b01001000101101: pixel[2:0] = 3'b000;
      14'b01001000101110: pixel[2:0] = 3'b000;
      14'b01001000101111: pixel[2:0] = 3'b000;
      14'b01001000110000: pixel[2:0] = 3'b000;
      14'b01001000110001: pixel[2:0] = 3'b000;
      14'b01001000110010: pixel[2:0] = 3'b111;
      14'b01001000110011: pixel[2:0] = 3'b111;
      14'b01001000110100: pixel[2:0] = 3'b111;
      14'b01001000110101: pixel[2:0] = 3'b111;
      14'b01001000110110: pixel[2:0] = 3'b000;
      14'b01001000110111: pixel[2:0] = 3'b000;
      14'b01001000111000: pixel[2:0] = 3'b000;
      14'b01001000111001: pixel[2:0] = 3'b111;
      14'b01001000111010: pixel[2:0] = 3'b111;
      14'b01001000111011: pixel[2:0] = 3'b111;
      14'b01001000111100: pixel[2:0] = 3'b111;
      14'b01001000111101: pixel[2:0] = 3'b000;
      14'b01001000111110: pixel[2:0] = 3'b000;
      14'b01001000111111: pixel[2:0] = 3'b000;
      14'b01001001000000: pixel[2:0] = 3'b000;
      14'b01001001000001: pixel[2:0] = 3'b000;
      14'b01001001000010: pixel[2:0] = 3'b000;
      14'b01001001000011: pixel[2:0] = 3'b000;
      14'b01001001000100: pixel[2:0] = 3'b000;
      14'b01001001000101: pixel[2:0] = 3'b000;
      14'b01001001000110: pixel[2:0] = 3'b111;
      14'b01001001000111: pixel[2:0] = 3'b111;
      14'b01001001001000: pixel[2:0] = 3'b111;
      14'b01001001001001: pixel[2:0] = 3'b111;
      14'b01001001001010: pixel[2:0] = 3'b111;
      14'b01001001001011: pixel[2:0] = 3'b000;
      14'b01001001001100: pixel[2:0] = 3'b111;
      14'b01001001001101: pixel[2:0] = 3'b111;
      14'b01001001001110: pixel[2:0] = 3'b111;
      14'b01001001001111: pixel[2:0] = 3'b111;
      14'b01001001010000: pixel[2:0] = 3'b000;
      14'b01001001010001: pixel[2:0] = 3'b000;
      14'b01001001010010: pixel[2:0] = 3'b000;
      14'b01001001010011: pixel[2:0] = 3'b000;
      14'b01001001010100: pixel[2:0] = 3'b000;
      14'b01001001010101: pixel[2:0] = 3'b000;
      14'b01001001010110: pixel[2:0] = 3'b000;
      14'b01001001010111: pixel[2:0] = 3'b000;
      14'b01001001011000: pixel[2:0] = 3'b000;
      14'b01001001011001: pixel[2:0] = 3'b000;
      14'b01001001011010: pixel[2:0] = 3'b111;
      14'b01001001011011: pixel[2:0] = 3'b111;
      14'b01001001011100: pixel[2:0] = 3'b111;
      14'b01001001011101: pixel[2:0] = 3'b111;
      14'b01001001011110: pixel[2:0] = 3'b111;
      14'b01001001011111: pixel[2:0] = 3'b000;
      14'b01001001100000: pixel[2:0] = 3'b000;
      14'b01001001100001: pixel[2:0] = 3'b000;
      14'b01001001100010: pixel[2:0] = 3'b000;
      14'b01001001100011: pixel[2:0] = 3'b000;
      14'b01001001100100: pixel[2:0] = 3'b000;
      14'b01001001100101: pixel[2:0] = 3'b000;
      14'b01001001100110: pixel[2:0] = 3'b000;
      14'b01001001100111: pixel[2:0] = 3'b000;
      14'b01001001101000: pixel[2:0] = 3'b000;
      14'b01001001101001: pixel[2:0] = 3'b000;
      14'b01001001101010: pixel[2:0] = 3'b000;
      14'b01001001101011: pixel[2:0] = 3'b000;
      14'b01001001101100: pixel[2:0] = 3'b000;
      14'b01001001101101: pixel[2:0] = 3'b000;
      14'b01001001101110: pixel[2:0] = 3'b000;
      14'b01001001101111: pixel[2:0] = 3'b000;
      14'b01001001110000: pixel[2:0] = 3'b111;
      14'b01001001110001: pixel[2:0] = 3'b111;
      14'b01001001110010: pixel[2:0] = 3'b111;
      14'b01001001110011: pixel[2:0] = 3'b111;
      14'b01001001110100: pixel[2:0] = 3'b111;
      14'b01001001110101: pixel[2:0] = 3'b000;
      14'b01001001110110: pixel[2:0] = 3'b000;
      14'b01001001110111: pixel[2:0] = 3'b000;
      14'b01001001111000: pixel[2:0] = 3'b000;
      14'b01001001111001: pixel[2:0] = 3'b000;
      14'b01001001111010: pixel[2:0] = 3'b000;
      14'b01001001111011: pixel[2:0] = 3'b000;
      14'b01001001111100: pixel[2:0] = 3'b000;
      14'b01001001111101: pixel[2:0] = 3'b111;
      14'b01001001111110: pixel[2:0] = 3'b111;
      14'b01001001111111: pixel[2:0] = 3'b111;
      14'b01001010000000: pixel[2:0] = 3'b111;
      14'b01001010000001: pixel[2:0] = 3'b111;
      14'b01001010000010: pixel[2:0] = 3'b111;
      14'b01001010000011: pixel[2:0] = 3'b000;
      14'b01001010000100: pixel[2:0] = 3'b000;
      14'b01001010000101: pixel[2:0] = 3'b000;
      14'b01001010000110: pixel[2:0] = 3'b000;
      14'b01001010000111: pixel[2:0] = 3'b000;
      14'b01001100000000: pixel[2:0] = 3'b000;
      14'b01001100000001: pixel[2:0] = 3'b000;
      14'b01001100000010: pixel[2:0] = 3'b111;
      14'b01001100000011: pixel[2:0] = 3'b111;
      14'b01001100000100: pixel[2:0] = 3'b111;
      14'b01001100000101: pixel[2:0] = 3'b111;
      14'b01001100000110: pixel[2:0] = 3'b111;
      14'b01001100000111: pixel[2:0] = 3'b000;
      14'b01001100001000: pixel[2:0] = 3'b000;
      14'b01001100001001: pixel[2:0] = 3'b000;
      14'b01001100001010: pixel[2:0] = 3'b000;
      14'b01001100001011: pixel[2:0] = 3'b000;
      14'b01001100001100: pixel[2:0] = 3'b000;
      14'b01001100001101: pixel[2:0] = 3'b000;
      14'b01001100001110: pixel[2:0] = 3'b000;
      14'b01001100001111: pixel[2:0] = 3'b111;
      14'b01001100010000: pixel[2:0] = 3'b111;
      14'b01001100010001: pixel[2:0] = 3'b111;
      14'b01001100010010: pixel[2:0] = 3'b111;
      14'b01001100010011: pixel[2:0] = 3'b111;
      14'b01001100010100: pixel[2:0] = 3'b000;
      14'b01001100010101: pixel[2:0] = 3'b000;
      14'b01001100010110: pixel[2:0] = 3'b000;
      14'b01001100010111: pixel[2:0] = 3'b000;
      14'b01001100011000: pixel[2:0] = 3'b000;
      14'b01001100011001: pixel[2:0] = 3'b111;
      14'b01001100011010: pixel[2:0] = 3'b111;
      14'b01001100011011: pixel[2:0] = 3'b111;
      14'b01001100011100: pixel[2:0] = 3'b111;
      14'b01001100011101: pixel[2:0] = 3'b111;
      14'b01001100011110: pixel[2:0] = 3'b000;
      14'b01001100011111: pixel[2:0] = 3'b000;
      14'b01001100100000: pixel[2:0] = 3'b000;
      14'b01001100100001: pixel[2:0] = 3'b000;
      14'b01001100100010: pixel[2:0] = 3'b000;
      14'b01001100100011: pixel[2:0] = 3'b000;
      14'b01001100100100: pixel[2:0] = 3'b000;
      14'b01001100100101: pixel[2:0] = 3'b000;
      14'b01001100100110: pixel[2:0] = 3'b000;
      14'b01001100100111: pixel[2:0] = 3'b000;
      14'b01001100101000: pixel[2:0] = 3'b000;
      14'b01001100101001: pixel[2:0] = 3'b000;
      14'b01001100101010: pixel[2:0] = 3'b000;
      14'b01001100101011: pixel[2:0] = 3'b000;
      14'b01001100101100: pixel[2:0] = 3'b000;
      14'b01001100101101: pixel[2:0] = 3'b000;
      14'b01001100101110: pixel[2:0] = 3'b000;
      14'b01001100101111: pixel[2:0] = 3'b000;
      14'b01001100110000: pixel[2:0] = 3'b000;
      14'b01001100110001: pixel[2:0] = 3'b000;
      14'b01001100110010: pixel[2:0] = 3'b111;
      14'b01001100110011: pixel[2:0] = 3'b111;
      14'b01001100110100: pixel[2:0] = 3'b111;
      14'b01001100110101: pixel[2:0] = 3'b111;
      14'b01001100110110: pixel[2:0] = 3'b000;
      14'b01001100110111: pixel[2:0] = 3'b000;
      14'b01001100111000: pixel[2:0] = 3'b000;
      14'b01001100111001: pixel[2:0] = 3'b111;
      14'b01001100111010: pixel[2:0] = 3'b111;
      14'b01001100111011: pixel[2:0] = 3'b111;
      14'b01001100111100: pixel[2:0] = 3'b111;
      14'b01001100111101: pixel[2:0] = 3'b111;
      14'b01001100111110: pixel[2:0] = 3'b000;
      14'b01001100111111: pixel[2:0] = 3'b000;
      14'b01001101000000: pixel[2:0] = 3'b000;
      14'b01001101000001: pixel[2:0] = 3'b000;
      14'b01001101000010: pixel[2:0] = 3'b000;
      14'b01001101000011: pixel[2:0] = 3'b000;
      14'b01001101000100: pixel[2:0] = 3'b000;
      14'b01001101000101: pixel[2:0] = 3'b000;
      14'b01001101000110: pixel[2:0] = 3'b000;
      14'b01001101000111: pixel[2:0] = 3'b111;
      14'b01001101001000: pixel[2:0] = 3'b111;
      14'b01001101001001: pixel[2:0] = 3'b111;
      14'b01001101001010: pixel[2:0] = 3'b111;
      14'b01001101001011: pixel[2:0] = 3'b111;
      14'b01001101001100: pixel[2:0] = 3'b111;
      14'b01001101001101: pixel[2:0] = 3'b111;
      14'b01001101001110: pixel[2:0] = 3'b111;
      14'b01001101001111: pixel[2:0] = 3'b111;
      14'b01001101010000: pixel[2:0] = 3'b000;
      14'b01001101010001: pixel[2:0] = 3'b000;
      14'b01001101010010: pixel[2:0] = 3'b000;
      14'b01001101010011: pixel[2:0] = 3'b000;
      14'b01001101010100: pixel[2:0] = 3'b000;
      14'b01001101010101: pixel[2:0] = 3'b000;
      14'b01001101010110: pixel[2:0] = 3'b000;
      14'b01001101010111: pixel[2:0] = 3'b000;
      14'b01001101011000: pixel[2:0] = 3'b000;
      14'b01001101011001: pixel[2:0] = 3'b000;
      14'b01001101011010: pixel[2:0] = 3'b111;
      14'b01001101011011: pixel[2:0] = 3'b111;
      14'b01001101011100: pixel[2:0] = 3'b111;
      14'b01001101011101: pixel[2:0] = 3'b111;
      14'b01001101011110: pixel[2:0] = 3'b111;
      14'b01001101011111: pixel[2:0] = 3'b111;
      14'b01001101100000: pixel[2:0] = 3'b111;
      14'b01001101100001: pixel[2:0] = 3'b111;
      14'b01001101100010: pixel[2:0] = 3'b111;
      14'b01001101100011: pixel[2:0] = 3'b111;
      14'b01001101100100: pixel[2:0] = 3'b111;
      14'b01001101100101: pixel[2:0] = 3'b111;
      14'b01001101100110: pixel[2:0] = 3'b111;
      14'b01001101100111: pixel[2:0] = 3'b111;
      14'b01001101101000: pixel[2:0] = 3'b111;
      14'b01001101101001: pixel[2:0] = 3'b000;
      14'b01001101101010: pixel[2:0] = 3'b000;
      14'b01001101101011: pixel[2:0] = 3'b000;
      14'b01001101101100: pixel[2:0] = 3'b000;
      14'b01001101101101: pixel[2:0] = 3'b000;
      14'b01001101101110: pixel[2:0] = 3'b000;
      14'b01001101101111: pixel[2:0] = 3'b000;
      14'b01001101110000: pixel[2:0] = 3'b111;
      14'b01001101110001: pixel[2:0] = 3'b111;
      14'b01001101110010: pixel[2:0] = 3'b111;
      14'b01001101110011: pixel[2:0] = 3'b111;
      14'b01001101110100: pixel[2:0] = 3'b111;
      14'b01001101110101: pixel[2:0] = 3'b000;
      14'b01001101110110: pixel[2:0] = 3'b000;
      14'b01001101110111: pixel[2:0] = 3'b000;
      14'b01001101111000: pixel[2:0] = 3'b000;
      14'b01001101111001: pixel[2:0] = 3'b000;
      14'b01001101111010: pixel[2:0] = 3'b000;
      14'b01001101111011: pixel[2:0] = 3'b000;
      14'b01001101111100: pixel[2:0] = 3'b000;
      14'b01001101111101: pixel[2:0] = 3'b111;
      14'b01001101111110: pixel[2:0] = 3'b111;
      14'b01001101111111: pixel[2:0] = 3'b111;
      14'b01001110000000: pixel[2:0] = 3'b111;
      14'b01001110000001: pixel[2:0] = 3'b111;
      14'b01001110000010: pixel[2:0] = 3'b000;
      14'b01001110000011: pixel[2:0] = 3'b000;
      14'b01001110000100: pixel[2:0] = 3'b000;
      14'b01001110000101: pixel[2:0] = 3'b000;
      14'b01001110000110: pixel[2:0] = 3'b000;
      14'b01001110000111: pixel[2:0] = 3'b000;
      14'b01010000000000: pixel[2:0] = 3'b000;
      14'b01010000000001: pixel[2:0] = 3'b000;
      14'b01010000000010: pixel[2:0] = 3'b111;
      14'b01010000000011: pixel[2:0] = 3'b111;
      14'b01010000000100: pixel[2:0] = 3'b111;
      14'b01010000000101: pixel[2:0] = 3'b111;
      14'b01010000000110: pixel[2:0] = 3'b111;
      14'b01010000000111: pixel[2:0] = 3'b000;
      14'b01010000001000: pixel[2:0] = 3'b000;
      14'b01010000001001: pixel[2:0] = 3'b000;
      14'b01010000001010: pixel[2:0] = 3'b000;
      14'b01010000001011: pixel[2:0] = 3'b000;
      14'b01010000001100: pixel[2:0] = 3'b000;
      14'b01010000001101: pixel[2:0] = 3'b000;
      14'b01010000001110: pixel[2:0] = 3'b111;
      14'b01010000001111: pixel[2:0] = 3'b111;
      14'b01010000010000: pixel[2:0] = 3'b111;
      14'b01010000010001: pixel[2:0] = 3'b111;
      14'b01010000010010: pixel[2:0] = 3'b111;
      14'b01010000010011: pixel[2:0] = 3'b111;
      14'b01010000010100: pixel[2:0] = 3'b000;
      14'b01010000010101: pixel[2:0] = 3'b000;
      14'b01010000010110: pixel[2:0] = 3'b000;
      14'b01010000010111: pixel[2:0] = 3'b000;
      14'b01010000011000: pixel[2:0] = 3'b000;
      14'b01010000011001: pixel[2:0] = 3'b111;
      14'b01010000011010: pixel[2:0] = 3'b111;
      14'b01010000011011: pixel[2:0] = 3'b111;
      14'b01010000011100: pixel[2:0] = 3'b111;
      14'b01010000011101: pixel[2:0] = 3'b111;
      14'b01010000011110: pixel[2:0] = 3'b000;
      14'b01010000011111: pixel[2:0] = 3'b000;
      14'b01010000100000: pixel[2:0] = 3'b000;
      14'b01010000100001: pixel[2:0] = 3'b000;
      14'b01010000100010: pixel[2:0] = 3'b000;
      14'b01010000100011: pixel[2:0] = 3'b000;
      14'b01010000100100: pixel[2:0] = 3'b000;
      14'b01010000100101: pixel[2:0] = 3'b000;
      14'b01010000100110: pixel[2:0] = 3'b000;
      14'b01010000100111: pixel[2:0] = 3'b000;
      14'b01010000101000: pixel[2:0] = 3'b000;
      14'b01010000101001: pixel[2:0] = 3'b000;
      14'b01010000101010: pixel[2:0] = 3'b000;
      14'b01010000101011: pixel[2:0] = 3'b000;
      14'b01010000101100: pixel[2:0] = 3'b000;
      14'b01010000101101: pixel[2:0] = 3'b000;
      14'b01010000101110: pixel[2:0] = 3'b000;
      14'b01010000101111: pixel[2:0] = 3'b000;
      14'b01010000110000: pixel[2:0] = 3'b000;
      14'b01010000110001: pixel[2:0] = 3'b000;
      14'b01010000110010: pixel[2:0] = 3'b111;
      14'b01010000110011: pixel[2:0] = 3'b111;
      14'b01010000110100: pixel[2:0] = 3'b111;
      14'b01010000110101: pixel[2:0] = 3'b111;
      14'b01010000110110: pixel[2:0] = 3'b000;
      14'b01010000110111: pixel[2:0] = 3'b000;
      14'b01010000111000: pixel[2:0] = 3'b000;
      14'b01010000111001: pixel[2:0] = 3'b000;
      14'b01010000111010: pixel[2:0] = 3'b111;
      14'b01010000111011: pixel[2:0] = 3'b111;
      14'b01010000111100: pixel[2:0] = 3'b111;
      14'b01010000111101: pixel[2:0] = 3'b111;
      14'b01010000111110: pixel[2:0] = 3'b000;
      14'b01010000111111: pixel[2:0] = 3'b000;
      14'b01010001000000: pixel[2:0] = 3'b000;
      14'b01010001000001: pixel[2:0] = 3'b000;
      14'b01010001000010: pixel[2:0] = 3'b000;
      14'b01010001000011: pixel[2:0] = 3'b000;
      14'b01010001000100: pixel[2:0] = 3'b000;
      14'b01010001000101: pixel[2:0] = 3'b000;
      14'b01010001000110: pixel[2:0] = 3'b000;
      14'b01010001000111: pixel[2:0] = 3'b111;
      14'b01010001001000: pixel[2:0] = 3'b111;
      14'b01010001001001: pixel[2:0] = 3'b111;
      14'b01010001001010: pixel[2:0] = 3'b111;
      14'b01010001001011: pixel[2:0] = 3'b111;
      14'b01010001001100: pixel[2:0] = 3'b111;
      14'b01010001001101: pixel[2:0] = 3'b111;
      14'b01010001001110: pixel[2:0] = 3'b111;
      14'b01010001001111: pixel[2:0] = 3'b000;
      14'b01010001010000: pixel[2:0] = 3'b000;
      14'b01010001010001: pixel[2:0] = 3'b000;
      14'b01010001010010: pixel[2:0] = 3'b000;
      14'b01010001010011: pixel[2:0] = 3'b000;
      14'b01010001010100: pixel[2:0] = 3'b000;
      14'b01010001010101: pixel[2:0] = 3'b000;
      14'b01010001010110: pixel[2:0] = 3'b000;
      14'b01010001010111: pixel[2:0] = 3'b000;
      14'b01010001011000: pixel[2:0] = 3'b000;
      14'b01010001011001: pixel[2:0] = 3'b000;
      14'b01010001011010: pixel[2:0] = 3'b111;
      14'b01010001011011: pixel[2:0] = 3'b111;
      14'b01010001011100: pixel[2:0] = 3'b111;
      14'b01010001011101: pixel[2:0] = 3'b111;
      14'b01010001011110: pixel[2:0] = 3'b111;
      14'b01010001011111: pixel[2:0] = 3'b111;
      14'b01010001100000: pixel[2:0] = 3'b111;
      14'b01010001100001: pixel[2:0] = 3'b111;
      14'b01010001100010: pixel[2:0] = 3'b111;
      14'b01010001100011: pixel[2:0] = 3'b111;
      14'b01010001100100: pixel[2:0] = 3'b111;
      14'b01010001100101: pixel[2:0] = 3'b111;
      14'b01010001100110: pixel[2:0] = 3'b111;
      14'b01010001100111: pixel[2:0] = 3'b111;
      14'b01010001101000: pixel[2:0] = 3'b111;
      14'b01010001101001: pixel[2:0] = 3'b000;
      14'b01010001101010: pixel[2:0] = 3'b000;
      14'b01010001101011: pixel[2:0] = 3'b000;
      14'b01010001101100: pixel[2:0] = 3'b000;
      14'b01010001101101: pixel[2:0] = 3'b000;
      14'b01010001101110: pixel[2:0] = 3'b000;
      14'b01010001101111: pixel[2:0] = 3'b000;
      14'b01010001110000: pixel[2:0] = 3'b111;
      14'b01010001110001: pixel[2:0] = 3'b111;
      14'b01010001110010: pixel[2:0] = 3'b111;
      14'b01010001110011: pixel[2:0] = 3'b111;
      14'b01010001110100: pixel[2:0] = 3'b111;
      14'b01010001110101: pixel[2:0] = 3'b111;
      14'b01010001110110: pixel[2:0] = 3'b111;
      14'b01010001110111: pixel[2:0] = 3'b111;
      14'b01010001111000: pixel[2:0] = 3'b111;
      14'b01010001111001: pixel[2:0] = 3'b111;
      14'b01010001111010: pixel[2:0] = 3'b111;
      14'b01010001111011: pixel[2:0] = 3'b111;
      14'b01010001111100: pixel[2:0] = 3'b111;
      14'b01010001111101: pixel[2:0] = 3'b111;
      14'b01010001111110: pixel[2:0] = 3'b111;
      14'b01010001111111: pixel[2:0] = 3'b111;
      14'b01010010000000: pixel[2:0] = 3'b111;
      14'b01010010000001: pixel[2:0] = 3'b111;
      14'b01010010000010: pixel[2:0] = 3'b000;
      14'b01010010000011: pixel[2:0] = 3'b000;
      14'b01010010000100: pixel[2:0] = 3'b000;
      14'b01010010000101: pixel[2:0] = 3'b000;
      14'b01010010000110: pixel[2:0] = 3'b000;
      14'b01010010000111: pixel[2:0] = 3'b000;
      14'b01010100000000: pixel[2:0] = 3'b000;
      14'b01010100000001: pixel[2:0] = 3'b000;
      14'b01010100000010: pixel[2:0] = 3'b111;
      14'b01010100000011: pixel[2:0] = 3'b111;
      14'b01010100000100: pixel[2:0] = 3'b111;
      14'b01010100000101: pixel[2:0] = 3'b111;
      14'b01010100000110: pixel[2:0] = 3'b111;
      14'b01010100000111: pixel[2:0] = 3'b111;
      14'b01010100001000: pixel[2:0] = 3'b111;
      14'b01010100001001: pixel[2:0] = 3'b111;
      14'b01010100001010: pixel[2:0] = 3'b111;
      14'b01010100001011: pixel[2:0] = 3'b111;
      14'b01010100001100: pixel[2:0] = 3'b111;
      14'b01010100001101: pixel[2:0] = 3'b111;
      14'b01010100001110: pixel[2:0] = 3'b111;
      14'b01010100001111: pixel[2:0] = 3'b111;
      14'b01010100010000: pixel[2:0] = 3'b111;
      14'b01010100010001: pixel[2:0] = 3'b111;
      14'b01010100010010: pixel[2:0] = 3'b111;
      14'b01010100010011: pixel[2:0] = 3'b000;
      14'b01010100010100: pixel[2:0] = 3'b000;
      14'b01010100010101: pixel[2:0] = 3'b000;
      14'b01010100010110: pixel[2:0] = 3'b000;
      14'b01010100010111: pixel[2:0] = 3'b000;
      14'b01010100011000: pixel[2:0] = 3'b000;
      14'b01010100011001: pixel[2:0] = 3'b111;
      14'b01010100011010: pixel[2:0] = 3'b111;
      14'b01010100011011: pixel[2:0] = 3'b111;
      14'b01010100011100: pixel[2:0] = 3'b111;
      14'b01010100011101: pixel[2:0] = 3'b111;
      14'b01010100011110: pixel[2:0] = 3'b000;
      14'b01010100011111: pixel[2:0] = 3'b000;
      14'b01010100100000: pixel[2:0] = 3'b000;
      14'b01010100100001: pixel[2:0] = 3'b000;
      14'b01010100100010: pixel[2:0] = 3'b000;
      14'b01010100100011: pixel[2:0] = 3'b000;
      14'b01010100100100: pixel[2:0] = 3'b000;
      14'b01010100100101: pixel[2:0] = 3'b000;
      14'b01010100100110: pixel[2:0] = 3'b000;
      14'b01010100100111: pixel[2:0] = 3'b000;
      14'b01010100101000: pixel[2:0] = 3'b000;
      14'b01010100101001: pixel[2:0] = 3'b000;
      14'b01010100101010: pixel[2:0] = 3'b000;
      14'b01010100101011: pixel[2:0] = 3'b000;
      14'b01010100101100: pixel[2:0] = 3'b000;
      14'b01010100101101: pixel[2:0] = 3'b000;
      14'b01010100101110: pixel[2:0] = 3'b000;
      14'b01010100101111: pixel[2:0] = 3'b000;
      14'b01010100110000: pixel[2:0] = 3'b000;
      14'b01010100110001: pixel[2:0] = 3'b111;
      14'b01010100110010: pixel[2:0] = 3'b111;
      14'b01010100110011: pixel[2:0] = 3'b111;
      14'b01010100110100: pixel[2:0] = 3'b111;
      14'b01010100110101: pixel[2:0] = 3'b111;
      14'b01010100110110: pixel[2:0] = 3'b000;
      14'b01010100110111: pixel[2:0] = 3'b000;
      14'b01010100111000: pixel[2:0] = 3'b000;
      14'b01010100111001: pixel[2:0] = 3'b000;
      14'b01010100111010: pixel[2:0] = 3'b111;
      14'b01010100111011: pixel[2:0] = 3'b111;
      14'b01010100111100: pixel[2:0] = 3'b111;
      14'b01010100111101: pixel[2:0] = 3'b111;
      14'b01010100111110: pixel[2:0] = 3'b000;
      14'b01010100111111: pixel[2:0] = 3'b000;
      14'b01010101000000: pixel[2:0] = 3'b000;
      14'b01010101000001: pixel[2:0] = 3'b000;
      14'b01010101000010: pixel[2:0] = 3'b000;
      14'b01010101000011: pixel[2:0] = 3'b000;
      14'b01010101000100: pixel[2:0] = 3'b000;
      14'b01010101000101: pixel[2:0] = 3'b000;
      14'b01010101000110: pixel[2:0] = 3'b000;
      14'b01010101000111: pixel[2:0] = 3'b111;
      14'b01010101001000: pixel[2:0] = 3'b111;
      14'b01010101001001: pixel[2:0] = 3'b111;
      14'b01010101001010: pixel[2:0] = 3'b111;
      14'b01010101001011: pixel[2:0] = 3'b111;
      14'b01010101001100: pixel[2:0] = 3'b111;
      14'b01010101001101: pixel[2:0] = 3'b111;
      14'b01010101001110: pixel[2:0] = 3'b111;
      14'b01010101001111: pixel[2:0] = 3'b000;
      14'b01010101010000: pixel[2:0] = 3'b000;
      14'b01010101010001: pixel[2:0] = 3'b000;
      14'b01010101010010: pixel[2:0] = 3'b000;
      14'b01010101010011: pixel[2:0] = 3'b000;
      14'b01010101010100: pixel[2:0] = 3'b000;
      14'b01010101010101: pixel[2:0] = 3'b000;
      14'b01010101010110: pixel[2:0] = 3'b000;
      14'b01010101010111: pixel[2:0] = 3'b000;
      14'b01010101011000: pixel[2:0] = 3'b000;
      14'b01010101011001: pixel[2:0] = 3'b000;
      14'b01010101011010: pixel[2:0] = 3'b111;
      14'b01010101011011: pixel[2:0] = 3'b111;
      14'b01010101011100: pixel[2:0] = 3'b111;
      14'b01010101011101: pixel[2:0] = 3'b111;
      14'b01010101011110: pixel[2:0] = 3'b111;
      14'b01010101011111: pixel[2:0] = 3'b111;
      14'b01010101100000: pixel[2:0] = 3'b111;
      14'b01010101100001: pixel[2:0] = 3'b111;
      14'b01010101100010: pixel[2:0] = 3'b111;
      14'b01010101100011: pixel[2:0] = 3'b111;
      14'b01010101100100: pixel[2:0] = 3'b111;
      14'b01010101100101: pixel[2:0] = 3'b111;
      14'b01010101100110: pixel[2:0] = 3'b111;
      14'b01010101100111: pixel[2:0] = 3'b111;
      14'b01010101101000: pixel[2:0] = 3'b111;
      14'b01010101101001: pixel[2:0] = 3'b000;
      14'b01010101101010: pixel[2:0] = 3'b000;
      14'b01010101101011: pixel[2:0] = 3'b000;
      14'b01010101101100: pixel[2:0] = 3'b000;
      14'b01010101101101: pixel[2:0] = 3'b000;
      14'b01010101101110: pixel[2:0] = 3'b000;
      14'b01010101101111: pixel[2:0] = 3'b000;
      14'b01010101110000: pixel[2:0] = 3'b111;
      14'b01010101110001: pixel[2:0] = 3'b111;
      14'b01010101110010: pixel[2:0] = 3'b111;
      14'b01010101110011: pixel[2:0] = 3'b111;
      14'b01010101110100: pixel[2:0] = 3'b111;
      14'b01010101110101: pixel[2:0] = 3'b111;
      14'b01010101110110: pixel[2:0] = 3'b111;
      14'b01010101110111: pixel[2:0] = 3'b111;
      14'b01010101111000: pixel[2:0] = 3'b111;
      14'b01010101111001: pixel[2:0] = 3'b111;
      14'b01010101111010: pixel[2:0] = 3'b111;
      14'b01010101111011: pixel[2:0] = 3'b111;
      14'b01010101111100: pixel[2:0] = 3'b111;
      14'b01010101111101: pixel[2:0] = 3'b111;
      14'b01010101111110: pixel[2:0] = 3'b111;
      14'b01010101111111: pixel[2:0] = 3'b111;
      14'b01010110000000: pixel[2:0] = 3'b111;
      14'b01010110000001: pixel[2:0] = 3'b000;
      14'b01010110000010: pixel[2:0] = 3'b000;
      14'b01010110000011: pixel[2:0] = 3'b000;
      14'b01010110000100: pixel[2:0] = 3'b000;
      14'b01010110000101: pixel[2:0] = 3'b000;
      14'b01010110000110: pixel[2:0] = 3'b000;
      14'b01010110000111: pixel[2:0] = 3'b000;
      14'b01011000000000: pixel[2:0] = 3'b000;
      14'b01011000000001: pixel[2:0] = 3'b000;
      14'b01011000000010: pixel[2:0] = 3'b111;
      14'b01011000000011: pixel[2:0] = 3'b111;
      14'b01011000000100: pixel[2:0] = 3'b111;
      14'b01011000000101: pixel[2:0] = 3'b111;
      14'b01011000000110: pixel[2:0] = 3'b111;
      14'b01011000000111: pixel[2:0] = 3'b111;
      14'b01011000001000: pixel[2:0] = 3'b111;
      14'b01011000001001: pixel[2:0] = 3'b111;
      14'b01011000001010: pixel[2:0] = 3'b111;
      14'b01011000001011: pixel[2:0] = 3'b111;
      14'b01011000001100: pixel[2:0] = 3'b111;
      14'b01011000001101: pixel[2:0] = 3'b111;
      14'b01011000001110: pixel[2:0] = 3'b111;
      14'b01011000001111: pixel[2:0] = 3'b111;
      14'b01011000010000: pixel[2:0] = 3'b111;
      14'b01011000010001: pixel[2:0] = 3'b111;
      14'b01011000010010: pixel[2:0] = 3'b111;
      14'b01011000010011: pixel[2:0] = 3'b000;
      14'b01011000010100: pixel[2:0] = 3'b000;
      14'b01011000010101: pixel[2:0] = 3'b000;
      14'b01011000010110: pixel[2:0] = 3'b000;
      14'b01011000010111: pixel[2:0] = 3'b000;
      14'b01011000011000: pixel[2:0] = 3'b000;
      14'b01011000011001: pixel[2:0] = 3'b111;
      14'b01011000011010: pixel[2:0] = 3'b111;
      14'b01011000011011: pixel[2:0] = 3'b111;
      14'b01011000011100: pixel[2:0] = 3'b111;
      14'b01011000011101: pixel[2:0] = 3'b111;
      14'b01011000011110: pixel[2:0] = 3'b000;
      14'b01011000011111: pixel[2:0] = 3'b000;
      14'b01011000100000: pixel[2:0] = 3'b000;
      14'b01011000100001: pixel[2:0] = 3'b000;
      14'b01011000100010: pixel[2:0] = 3'b000;
      14'b01011000100011: pixel[2:0] = 3'b000;
      14'b01011000100100: pixel[2:0] = 3'b000;
      14'b01011000100101: pixel[2:0] = 3'b000;
      14'b01011000100110: pixel[2:0] = 3'b000;
      14'b01011000100111: pixel[2:0] = 3'b000;
      14'b01011000101000: pixel[2:0] = 3'b000;
      14'b01011000101001: pixel[2:0] = 3'b000;
      14'b01011000101010: pixel[2:0] = 3'b000;
      14'b01011000101011: pixel[2:0] = 3'b000;
      14'b01011000101100: pixel[2:0] = 3'b000;
      14'b01011000101101: pixel[2:0] = 3'b000;
      14'b01011000101110: pixel[2:0] = 3'b000;
      14'b01011000101111: pixel[2:0] = 3'b000;
      14'b01011000110000: pixel[2:0] = 3'b000;
      14'b01011000110001: pixel[2:0] = 3'b111;
      14'b01011000110010: pixel[2:0] = 3'b111;
      14'b01011000110011: pixel[2:0] = 3'b111;
      14'b01011000110100: pixel[2:0] = 3'b111;
      14'b01011000110101: pixel[2:0] = 3'b000;
      14'b01011000110110: pixel[2:0] = 3'b000;
      14'b01011000110111: pixel[2:0] = 3'b000;
      14'b01011000111000: pixel[2:0] = 3'b000;
      14'b01011000111001: pixel[2:0] = 3'b000;
      14'b01011000111010: pixel[2:0] = 3'b111;
      14'b01011000111011: pixel[2:0] = 3'b111;
      14'b01011000111100: pixel[2:0] = 3'b111;
      14'b01011000111101: pixel[2:0] = 3'b111;
      14'b01011000111110: pixel[2:0] = 3'b000;
      14'b01011000111111: pixel[2:0] = 3'b000;
      14'b01011001000000: pixel[2:0] = 3'b000;
      14'b01011001000001: pixel[2:0] = 3'b000;
      14'b01011001000010: pixel[2:0] = 3'b000;
      14'b01011001000011: pixel[2:0] = 3'b000;
      14'b01011001000100: pixel[2:0] = 3'b000;
      14'b01011001000101: pixel[2:0] = 3'b000;
      14'b01011001000110: pixel[2:0] = 3'b000;
      14'b01011001000111: pixel[2:0] = 3'b000;
      14'b01011001001000: pixel[2:0] = 3'b111;
      14'b01011001001001: pixel[2:0] = 3'b111;
      14'b01011001001010: pixel[2:0] = 3'b111;
      14'b01011001001011: pixel[2:0] = 3'b111;
      14'b01011001001100: pixel[2:0] = 3'b111;
      14'b01011001001101: pixel[2:0] = 3'b111;
      14'b01011001001110: pixel[2:0] = 3'b111;
      14'b01011001001111: pixel[2:0] = 3'b000;
      14'b01011001010000: pixel[2:0] = 3'b000;
      14'b01011001010001: pixel[2:0] = 3'b000;
      14'b01011001010010: pixel[2:0] = 3'b000;
      14'b01011001010011: pixel[2:0] = 3'b000;
      14'b01011001010100: pixel[2:0] = 3'b000;
      14'b01011001010101: pixel[2:0] = 3'b000;
      14'b01011001010110: pixel[2:0] = 3'b000;
      14'b01011001010111: pixel[2:0] = 3'b000;
      14'b01011001011000: pixel[2:0] = 3'b000;
      14'b01011001011001: pixel[2:0] = 3'b000;
      14'b01011001011010: pixel[2:0] = 3'b111;
      14'b01011001011011: pixel[2:0] = 3'b111;
      14'b01011001011100: pixel[2:0] = 3'b111;
      14'b01011001011101: pixel[2:0] = 3'b111;
      14'b01011001011110: pixel[2:0] = 3'b111;
      14'b01011001011111: pixel[2:0] = 3'b111;
      14'b01011001100000: pixel[2:0] = 3'b111;
      14'b01011001100001: pixel[2:0] = 3'b111;
      14'b01011001100010: pixel[2:0] = 3'b111;
      14'b01011001100011: pixel[2:0] = 3'b111;
      14'b01011001100100: pixel[2:0] = 3'b111;
      14'b01011001100101: pixel[2:0] = 3'b111;
      14'b01011001100110: pixel[2:0] = 3'b111;
      14'b01011001100111: pixel[2:0] = 3'b111;
      14'b01011001101000: pixel[2:0] = 3'b111;
      14'b01011001101001: pixel[2:0] = 3'b000;
      14'b01011001101010: pixel[2:0] = 3'b000;
      14'b01011001101011: pixel[2:0] = 3'b000;
      14'b01011001101100: pixel[2:0] = 3'b000;
      14'b01011001101101: pixel[2:0] = 3'b000;
      14'b01011001101110: pixel[2:0] = 3'b000;
      14'b01011001101111: pixel[2:0] = 3'b000;
      14'b01011001110000: pixel[2:0] = 3'b111;
      14'b01011001110001: pixel[2:0] = 3'b111;
      14'b01011001110010: pixel[2:0] = 3'b111;
      14'b01011001110011: pixel[2:0] = 3'b111;
      14'b01011001110100: pixel[2:0] = 3'b111;
      14'b01011001110101: pixel[2:0] = 3'b111;
      14'b01011001110110: pixel[2:0] = 3'b111;
      14'b01011001110111: pixel[2:0] = 3'b111;
      14'b01011001111000: pixel[2:0] = 3'b111;
      14'b01011001111001: pixel[2:0] = 3'b111;
      14'b01011001111010: pixel[2:0] = 3'b111;
      14'b01011001111011: pixel[2:0] = 3'b111;
      14'b01011001111100: pixel[2:0] = 3'b111;
      14'b01011001111101: pixel[2:0] = 3'b111;
      14'b01011001111110: pixel[2:0] = 3'b111;
      14'b01011001111111: pixel[2:0] = 3'b111;
      14'b01011010000000: pixel[2:0] = 3'b000;
      14'b01011010000001: pixel[2:0] = 3'b000;
      14'b01011010000010: pixel[2:0] = 3'b000;
      14'b01011010000011: pixel[2:0] = 3'b000;
      14'b01011010000100: pixel[2:0] = 3'b000;
      14'b01011010000101: pixel[2:0] = 3'b000;
      14'b01011010000110: pixel[2:0] = 3'b000;
      14'b01011010000111: pixel[2:0] = 3'b000;
      14'b01011100000000: pixel[2:0] = 3'b000;
      14'b01011100000001: pixel[2:0] = 3'b000;
      14'b01011100000010: pixel[2:0] = 3'b111;
      14'b01011100000011: pixel[2:0] = 3'b111;
      14'b01011100000100: pixel[2:0] = 3'b111;
      14'b01011100000101: pixel[2:0] = 3'b111;
      14'b01011100000110: pixel[2:0] = 3'b111;
      14'b01011100000111: pixel[2:0] = 3'b111;
      14'b01011100001000: pixel[2:0] = 3'b111;
      14'b01011100001001: pixel[2:0] = 3'b111;
      14'b01011100001010: pixel[2:0] = 3'b111;
      14'b01011100001011: pixel[2:0] = 3'b111;
      14'b01011100001100: pixel[2:0] = 3'b111;
      14'b01011100001101: pixel[2:0] = 3'b111;
      14'b01011100001110: pixel[2:0] = 3'b111;
      14'b01011100001111: pixel[2:0] = 3'b111;
      14'b01011100010000: pixel[2:0] = 3'b111;
      14'b01011100010001: pixel[2:0] = 3'b111;
      14'b01011100010010: pixel[2:0] = 3'b000;
      14'b01011100010011: pixel[2:0] = 3'b000;
      14'b01011100010100: pixel[2:0] = 3'b000;
      14'b01011100010101: pixel[2:0] = 3'b000;
      14'b01011100010110: pixel[2:0] = 3'b000;
      14'b01011100010111: pixel[2:0] = 3'b000;
      14'b01011100011000: pixel[2:0] = 3'b000;
      14'b01011100011001: pixel[2:0] = 3'b111;
      14'b01011100011010: pixel[2:0] = 3'b111;
      14'b01011100011011: pixel[2:0] = 3'b111;
      14'b01011100011100: pixel[2:0] = 3'b111;
      14'b01011100011101: pixel[2:0] = 3'b111;
      14'b01011100011110: pixel[2:0] = 3'b000;
      14'b01011100011111: pixel[2:0] = 3'b000;
      14'b01011100100000: pixel[2:0] = 3'b000;
      14'b01011100100001: pixel[2:0] = 3'b000;
      14'b01011100100010: pixel[2:0] = 3'b000;
      14'b01011100100011: pixel[2:0] = 3'b000;
      14'b01011100100100: pixel[2:0] = 3'b000;
      14'b01011100100101: pixel[2:0] = 3'b000;
      14'b01011100100110: pixel[2:0] = 3'b000;
      14'b01011100100111: pixel[2:0] = 3'b000;
      14'b01011100101000: pixel[2:0] = 3'b000;
      14'b01011100101001: pixel[2:0] = 3'b000;
      14'b01011100101010: pixel[2:0] = 3'b000;
      14'b01011100101011: pixel[2:0] = 3'b000;
      14'b01011100101100: pixel[2:0] = 3'b000;
      14'b01011100101101: pixel[2:0] = 3'b000;
      14'b01011100101110: pixel[2:0] = 3'b000;
      14'b01011100101111: pixel[2:0] = 3'b000;
      14'b01011100110000: pixel[2:0] = 3'b000;
      14'b01011100110001: pixel[2:0] = 3'b111;
      14'b01011100110010: pixel[2:0] = 3'b111;
      14'b01011100110011: pixel[2:0] = 3'b111;
      14'b01011100110100: pixel[2:0] = 3'b111;
      14'b01011100110101: pixel[2:0] = 3'b000;
      14'b01011100110110: pixel[2:0] = 3'b000;
      14'b01011100110111: pixel[2:0] = 3'b000;
      14'b01011100111000: pixel[2:0] = 3'b000;
      14'b01011100111001: pixel[2:0] = 3'b000;
      14'b01011100111010: pixel[2:0] = 3'b111;
      14'b01011100111011: pixel[2:0] = 3'b111;
      14'b01011100111100: pixel[2:0] = 3'b111;
      14'b01011100111101: pixel[2:0] = 3'b111;
      14'b01011100111110: pixel[2:0] = 3'b111;
      14'b01011100111111: pixel[2:0] = 3'b000;
      14'b01011101000000: pixel[2:0] = 3'b000;
      14'b01011101000001: pixel[2:0] = 3'b000;
      14'b01011101000010: pixel[2:0] = 3'b000;
      14'b01011101000011: pixel[2:0] = 3'b000;
      14'b01011101000100: pixel[2:0] = 3'b000;
      14'b01011101000101: pixel[2:0] = 3'b000;
      14'b01011101000110: pixel[2:0] = 3'b000;
      14'b01011101000111: pixel[2:0] = 3'b000;
      14'b01011101001000: pixel[2:0] = 3'b111;
      14'b01011101001001: pixel[2:0] = 3'b111;
      14'b01011101001010: pixel[2:0] = 3'b111;
      14'b01011101001011: pixel[2:0] = 3'b111;
      14'b01011101001100: pixel[2:0] = 3'b111;
      14'b01011101001101: pixel[2:0] = 3'b111;
      14'b01011101001110: pixel[2:0] = 3'b000;
      14'b01011101001111: pixel[2:0] = 3'b000;
      14'b01011101010000: pixel[2:0] = 3'b000;
      14'b01011101010001: pixel[2:0] = 3'b000;
      14'b01011101010010: pixel[2:0] = 3'b000;
      14'b01011101010011: pixel[2:0] = 3'b000;
      14'b01011101010100: pixel[2:0] = 3'b000;
      14'b01011101010101: pixel[2:0] = 3'b000;
      14'b01011101010110: pixel[2:0] = 3'b000;
      14'b01011101010111: pixel[2:0] = 3'b000;
      14'b01011101011000: pixel[2:0] = 3'b000;
      14'b01011101011001: pixel[2:0] = 3'b000;
      14'b01011101011010: pixel[2:0] = 3'b111;
      14'b01011101011011: pixel[2:0] = 3'b111;
      14'b01011101011100: pixel[2:0] = 3'b111;
      14'b01011101011101: pixel[2:0] = 3'b111;
      14'b01011101011110: pixel[2:0] = 3'b111;
      14'b01011101011111: pixel[2:0] = 3'b111;
      14'b01011101100000: pixel[2:0] = 3'b111;
      14'b01011101100001: pixel[2:0] = 3'b111;
      14'b01011101100010: pixel[2:0] = 3'b111;
      14'b01011101100011: pixel[2:0] = 3'b111;
      14'b01011101100100: pixel[2:0] = 3'b111;
      14'b01011101100101: pixel[2:0] = 3'b111;
      14'b01011101100110: pixel[2:0] = 3'b111;
      14'b01011101100111: pixel[2:0] = 3'b111;
      14'b01011101101000: pixel[2:0] = 3'b111;
      14'b01011101101001: pixel[2:0] = 3'b000;
      14'b01011101101010: pixel[2:0] = 3'b000;
      14'b01011101101011: pixel[2:0] = 3'b000;
      14'b01011101101100: pixel[2:0] = 3'b000;
      14'b01011101101101: pixel[2:0] = 3'b000;
      14'b01011101101110: pixel[2:0] = 3'b000;
      14'b01011101101111: pixel[2:0] = 3'b000;
      14'b01011101110000: pixel[2:0] = 3'b111;
      14'b01011101110001: pixel[2:0] = 3'b111;
      14'b01011101110010: pixel[2:0] = 3'b111;
      14'b01011101110011: pixel[2:0] = 3'b111;
      14'b01011101110100: pixel[2:0] = 3'b111;
      14'b01011101110101: pixel[2:0] = 3'b111;
      14'b01011101110110: pixel[2:0] = 3'b111;
      14'b01011101110111: pixel[2:0] = 3'b111;
      14'b01011101111000: pixel[2:0] = 3'b111;
      14'b01011101111001: pixel[2:0] = 3'b111;
      14'b01011101111010: pixel[2:0] = 3'b111;
      14'b01011101111011: pixel[2:0] = 3'b111;
      14'b01011101111100: pixel[2:0] = 3'b111;
      14'b01011101111101: pixel[2:0] = 3'b111;
      14'b01011101111110: pixel[2:0] = 3'b111;
      14'b01011101111111: pixel[2:0] = 3'b000;
      14'b01011110000000: pixel[2:0] = 3'b000;
      14'b01011110000001: pixel[2:0] = 3'b000;
      14'b01011110000010: pixel[2:0] = 3'b000;
      14'b01011110000011: pixel[2:0] = 3'b000;
      14'b01011110000100: pixel[2:0] = 3'b000;
      14'b01011110000101: pixel[2:0] = 3'b000;
      14'b01011110000110: pixel[2:0] = 3'b000;
      14'b01011110000111: pixel[2:0] = 3'b000;
      14'b01100000000000: pixel[2:0] = 3'b000;
      14'b01100000000001: pixel[2:0] = 3'b000;
      14'b01100000000010: pixel[2:0] = 3'b111;
      14'b01100000000011: pixel[2:0] = 3'b111;
      14'b01100000000100: pixel[2:0] = 3'b111;
      14'b01100000000101: pixel[2:0] = 3'b111;
      14'b01100000000110: pixel[2:0] = 3'b111;
      14'b01100000000111: pixel[2:0] = 3'b111;
      14'b01100000001000: pixel[2:0] = 3'b111;
      14'b01100000001001: pixel[2:0] = 3'b111;
      14'b01100000001010: pixel[2:0] = 3'b111;
      14'b01100000001011: pixel[2:0] = 3'b111;
      14'b01100000001100: pixel[2:0] = 3'b111;
      14'b01100000001101: pixel[2:0] = 3'b111;
      14'b01100000001110: pixel[2:0] = 3'b111;
      14'b01100000001111: pixel[2:0] = 3'b111;
      14'b01100000010000: pixel[2:0] = 3'b111;
      14'b01100000010001: pixel[2:0] = 3'b000;
      14'b01100000010010: pixel[2:0] = 3'b000;
      14'b01100000010011: pixel[2:0] = 3'b000;
      14'b01100000010100: pixel[2:0] = 3'b000;
      14'b01100000010101: pixel[2:0] = 3'b000;
      14'b01100000010110: pixel[2:0] = 3'b000;
      14'b01100000010111: pixel[2:0] = 3'b000;
      14'b01100000011000: pixel[2:0] = 3'b000;
      14'b01100000011001: pixel[2:0] = 3'b111;
      14'b01100000011010: pixel[2:0] = 3'b111;
      14'b01100000011011: pixel[2:0] = 3'b111;
      14'b01100000011100: pixel[2:0] = 3'b111;
      14'b01100000011101: pixel[2:0] = 3'b111;
      14'b01100000011110: pixel[2:0] = 3'b000;
      14'b01100000011111: pixel[2:0] = 3'b000;
      14'b01100000100000: pixel[2:0] = 3'b000;
      14'b01100000100001: pixel[2:0] = 3'b000;
      14'b01100000100010: pixel[2:0] = 3'b000;
      14'b01100000100011: pixel[2:0] = 3'b000;
      14'b01100000100100: pixel[2:0] = 3'b000;
      14'b01100000100101: pixel[2:0] = 3'b000;
      14'b01100000100110: pixel[2:0] = 3'b000;
      14'b01100000100111: pixel[2:0] = 3'b000;
      14'b01100000101000: pixel[2:0] = 3'b000;
      14'b01100000101001: pixel[2:0] = 3'b000;
      14'b01100000101010: pixel[2:0] = 3'b000;
      14'b01100000101011: pixel[2:0] = 3'b000;
      14'b01100000101100: pixel[2:0] = 3'b000;
      14'b01100000101101: pixel[2:0] = 3'b000;
      14'b01100000101110: pixel[2:0] = 3'b000;
      14'b01100000101111: pixel[2:0] = 3'b000;
      14'b01100000110000: pixel[2:0] = 3'b000;
      14'b01100000110001: pixel[2:0] = 3'b111;
      14'b01100000110010: pixel[2:0] = 3'b111;
      14'b01100000110011: pixel[2:0] = 3'b111;
      14'b01100000110100: pixel[2:0] = 3'b111;
      14'b01100000110101: pixel[2:0] = 3'b000;
      14'b01100000110110: pixel[2:0] = 3'b000;
      14'b01100000110111: pixel[2:0] = 3'b000;
      14'b01100000111000: pixel[2:0] = 3'b000;
      14'b01100000111001: pixel[2:0] = 3'b000;
      14'b01100000111010: pixel[2:0] = 3'b000;
      14'b01100000111011: pixel[2:0] = 3'b111;
      14'b01100000111100: pixel[2:0] = 3'b111;
      14'b01100000111101: pixel[2:0] = 3'b111;
      14'b01100000111110: pixel[2:0] = 3'b111;
      14'b01100000111111: pixel[2:0] = 3'b000;
      14'b01100001000000: pixel[2:0] = 3'b000;
      14'b01100001000001: pixel[2:0] = 3'b000;
      14'b01100001000010: pixel[2:0] = 3'b000;
      14'b01100001000011: pixel[2:0] = 3'b000;
      14'b01100001000100: pixel[2:0] = 3'b000;
      14'b01100001000101: pixel[2:0] = 3'b000;
      14'b01100001000110: pixel[2:0] = 3'b000;
      14'b01100001000111: pixel[2:0] = 3'b000;
      14'b01100001001000: pixel[2:0] = 3'b111;
      14'b01100001001001: pixel[2:0] = 3'b111;
      14'b01100001001010: pixel[2:0] = 3'b111;
      14'b01100001001011: pixel[2:0] = 3'b111;
      14'b01100001001100: pixel[2:0] = 3'b111;
      14'b01100001001101: pixel[2:0] = 3'b111;
      14'b01100001001110: pixel[2:0] = 3'b000;
      14'b01100001001111: pixel[2:0] = 3'b000;
      14'b01100001010000: pixel[2:0] = 3'b000;
      14'b01100001010001: pixel[2:0] = 3'b000;
      14'b01100001010010: pixel[2:0] = 3'b000;
      14'b01100001010011: pixel[2:0] = 3'b000;
      14'b01100001010100: pixel[2:0] = 3'b000;
      14'b01100001010101: pixel[2:0] = 3'b000;
      14'b01100001010110: pixel[2:0] = 3'b000;
      14'b01100001010111: pixel[2:0] = 3'b000;
      14'b01100001011000: pixel[2:0] = 3'b000;
      14'b01100001011001: pixel[2:0] = 3'b000;
      14'b01100001011010: pixel[2:0] = 3'b111;
      14'b01100001011011: pixel[2:0] = 3'b111;
      14'b01100001011100: pixel[2:0] = 3'b111;
      14'b01100001011101: pixel[2:0] = 3'b111;
      14'b01100001011110: pixel[2:0] = 3'b111;
      14'b01100001011111: pixel[2:0] = 3'b111;
      14'b01100001100000: pixel[2:0] = 3'b111;
      14'b01100001100001: pixel[2:0] = 3'b111;
      14'b01100001100010: pixel[2:0] = 3'b111;
      14'b01100001100011: pixel[2:0] = 3'b111;
      14'b01100001100100: pixel[2:0] = 3'b111;
      14'b01100001100101: pixel[2:0] = 3'b111;
      14'b01100001100110: pixel[2:0] = 3'b111;
      14'b01100001100111: pixel[2:0] = 3'b111;
      14'b01100001101000: pixel[2:0] = 3'b111;
      14'b01100001101001: pixel[2:0] = 3'b000;
      14'b01100001101010: pixel[2:0] = 3'b000;
      14'b01100001101011: pixel[2:0] = 3'b000;
      14'b01100001101100: pixel[2:0] = 3'b000;
      14'b01100001101101: pixel[2:0] = 3'b000;
      14'b01100001101110: pixel[2:0] = 3'b000;
      14'b01100001101111: pixel[2:0] = 3'b000;
      14'b01100001110000: pixel[2:0] = 3'b111;
      14'b01100001110001: pixel[2:0] = 3'b111;
      14'b01100001110010: pixel[2:0] = 3'b111;
      14'b01100001110011: pixel[2:0] = 3'b111;
      14'b01100001110100: pixel[2:0] = 3'b111;
      14'b01100001110101: pixel[2:0] = 3'b111;
      14'b01100001110110: pixel[2:0] = 3'b111;
      14'b01100001110111: pixel[2:0] = 3'b111;
      14'b01100001111000: pixel[2:0] = 3'b111;
      14'b01100001111001: pixel[2:0] = 3'b111;
      14'b01100001111010: pixel[2:0] = 3'b111;
      14'b01100001111011: pixel[2:0] = 3'b111;
      14'b01100001111100: pixel[2:0] = 3'b111;
      14'b01100001111101: pixel[2:0] = 3'b111;
      14'b01100001111110: pixel[2:0] = 3'b000;
      14'b01100001111111: pixel[2:0] = 3'b000;
      14'b01100010000000: pixel[2:0] = 3'b000;
      14'b01100010000001: pixel[2:0] = 3'b000;
      14'b01100010000010: pixel[2:0] = 3'b000;
      14'b01100010000011: pixel[2:0] = 3'b000;
      14'b01100010000100: pixel[2:0] = 3'b000;
      14'b01100010000101: pixel[2:0] = 3'b000;
      14'b01100010000110: pixel[2:0] = 3'b000;
      14'b01100010000111: pixel[2:0] = 3'b000;
      14'b01100100000000: pixel[2:0] = 3'b000;
      14'b01100100000001: pixel[2:0] = 3'b000;
      14'b01100100000010: pixel[2:0] = 3'b111;
      14'b01100100000011: pixel[2:0] = 3'b111;
      14'b01100100000100: pixel[2:0] = 3'b111;
      14'b01100100000101: pixel[2:0] = 3'b111;
      14'b01100100000110: pixel[2:0] = 3'b111;
      14'b01100100000111: pixel[2:0] = 3'b111;
      14'b01100100001000: pixel[2:0] = 3'b111;
      14'b01100100001001: pixel[2:0] = 3'b111;
      14'b01100100001010: pixel[2:0] = 3'b111;
      14'b01100100001011: pixel[2:0] = 3'b111;
      14'b01100100001100: pixel[2:0] = 3'b111;
      14'b01100100001101: pixel[2:0] = 3'b111;
      14'b01100100001110: pixel[2:0] = 3'b111;
      14'b01100100001111: pixel[2:0] = 3'b111;
      14'b01100100010000: pixel[2:0] = 3'b000;
      14'b01100100010001: pixel[2:0] = 3'b000;
      14'b01100100010010: pixel[2:0] = 3'b000;
      14'b01100100010011: pixel[2:0] = 3'b000;
      14'b01100100010100: pixel[2:0] = 3'b000;
      14'b01100100010101: pixel[2:0] = 3'b000;
      14'b01100100010110: pixel[2:0] = 3'b000;
      14'b01100100010111: pixel[2:0] = 3'b000;
      14'b01100100011000: pixel[2:0] = 3'b000;
      14'b01100100011001: pixel[2:0] = 3'b111;
      14'b01100100011010: pixel[2:0] = 3'b111;
      14'b01100100011011: pixel[2:0] = 3'b111;
      14'b01100100011100: pixel[2:0] = 3'b111;
      14'b01100100011101: pixel[2:0] = 3'b111;
      14'b01100100011110: pixel[2:0] = 3'b000;
      14'b01100100011111: pixel[2:0] = 3'b000;
      14'b01100100100000: pixel[2:0] = 3'b000;
      14'b01100100100001: pixel[2:0] = 3'b000;
      14'b01100100100010: pixel[2:0] = 3'b000;
      14'b01100100100011: pixel[2:0] = 3'b000;
      14'b01100100100100: pixel[2:0] = 3'b000;
      14'b01100100100101: pixel[2:0] = 3'b000;
      14'b01100100100110: pixel[2:0] = 3'b000;
      14'b01100100100111: pixel[2:0] = 3'b000;
      14'b01100100101000: pixel[2:0] = 3'b000;
      14'b01100100101001: pixel[2:0] = 3'b000;
      14'b01100100101010: pixel[2:0] = 3'b000;
      14'b01100100101011: pixel[2:0] = 3'b000;
      14'b01100100101100: pixel[2:0] = 3'b000;
      14'b01100100101101: pixel[2:0] = 3'b000;
      14'b01100100101110: pixel[2:0] = 3'b000;
      14'b01100100101111: pixel[2:0] = 3'b000;
      14'b01100100110000: pixel[2:0] = 3'b000;
      14'b01100100110001: pixel[2:0] = 3'b111;
      14'b01100100110010: pixel[2:0] = 3'b111;
      14'b01100100110011: pixel[2:0] = 3'b111;
      14'b01100100110100: pixel[2:0] = 3'b111;
      14'b01100100110101: pixel[2:0] = 3'b000;
      14'b01100100110110: pixel[2:0] = 3'b000;
      14'b01100100110111: pixel[2:0] = 3'b000;
      14'b01100100111000: pixel[2:0] = 3'b000;
      14'b01100100111001: pixel[2:0] = 3'b000;
      14'b01100100111010: pixel[2:0] = 3'b000;
      14'b01100100111011: pixel[2:0] = 3'b111;
      14'b01100100111100: pixel[2:0] = 3'b111;
      14'b01100100111101: pixel[2:0] = 3'b111;
      14'b01100100111110: pixel[2:0] = 3'b111;
      14'b01100100111111: pixel[2:0] = 3'b000;
      14'b01100101000000: pixel[2:0] = 3'b000;
      14'b01100101000001: pixel[2:0] = 3'b000;
      14'b01100101000010: pixel[2:0] = 3'b000;
      14'b01100101000011: pixel[2:0] = 3'b000;
      14'b01100101000100: pixel[2:0] = 3'b000;
      14'b01100101000101: pixel[2:0] = 3'b000;
      14'b01100101000110: pixel[2:0] = 3'b000;
      14'b01100101000111: pixel[2:0] = 3'b000;
      14'b01100101001000: pixel[2:0] = 3'b000;
      14'b01100101001001: pixel[2:0] = 3'b111;
      14'b01100101001010: pixel[2:0] = 3'b111;
      14'b01100101001011: pixel[2:0] = 3'b111;
      14'b01100101001100: pixel[2:0] = 3'b111;
      14'b01100101001101: pixel[2:0] = 3'b111;
      14'b01100101001110: pixel[2:0] = 3'b000;
      14'b01100101001111: pixel[2:0] = 3'b000;
      14'b01100101010000: pixel[2:0] = 3'b000;
      14'b01100101010001: pixel[2:0] = 3'b000;
      14'b01100101010010: pixel[2:0] = 3'b000;
      14'b01100101010011: pixel[2:0] = 3'b000;
      14'b01100101010100: pixel[2:0] = 3'b000;
      14'b01100101010101: pixel[2:0] = 3'b000;
      14'b01100101010110: pixel[2:0] = 3'b000;
      14'b01100101010111: pixel[2:0] = 3'b000;
      14'b01100101011000: pixel[2:0] = 3'b000;
      14'b01100101011001: pixel[2:0] = 3'b000;
      14'b01100101011010: pixel[2:0] = 3'b111;
      14'b01100101011011: pixel[2:0] = 3'b111;
      14'b01100101011100: pixel[2:0] = 3'b111;
      14'b01100101011101: pixel[2:0] = 3'b111;
      14'b01100101011110: pixel[2:0] = 3'b111;
      14'b01100101011111: pixel[2:0] = 3'b000;
      14'b01100101100000: pixel[2:0] = 3'b000;
      14'b01100101100001: pixel[2:0] = 3'b000;
      14'b01100101100010: pixel[2:0] = 3'b000;
      14'b01100101100011: pixel[2:0] = 3'b000;
      14'b01100101100100: pixel[2:0] = 3'b000;
      14'b01100101100101: pixel[2:0] = 3'b000;
      14'b01100101100110: pixel[2:0] = 3'b000;
      14'b01100101100111: pixel[2:0] = 3'b000;
      14'b01100101101000: pixel[2:0] = 3'b000;
      14'b01100101101001: pixel[2:0] = 3'b000;
      14'b01100101101010: pixel[2:0] = 3'b000;
      14'b01100101101011: pixel[2:0] = 3'b000;
      14'b01100101101100: pixel[2:0] = 3'b000;
      14'b01100101101101: pixel[2:0] = 3'b000;
      14'b01100101101110: pixel[2:0] = 3'b000;
      14'b01100101101111: pixel[2:0] = 3'b000;
      14'b01100101110000: pixel[2:0] = 3'b111;
      14'b01100101110001: pixel[2:0] = 3'b111;
      14'b01100101110010: pixel[2:0] = 3'b111;
      14'b01100101110011: pixel[2:0] = 3'b111;
      14'b01100101110100: pixel[2:0] = 3'b111;
      14'b01100101110101: pixel[2:0] = 3'b111;
      14'b01100101110110: pixel[2:0] = 3'b111;
      14'b01100101110111: pixel[2:0] = 3'b111;
      14'b01100101111000: pixel[2:0] = 3'b111;
      14'b01100101111001: pixel[2:0] = 3'b111;
      14'b01100101111010: pixel[2:0] = 3'b111;
      14'b01100101111011: pixel[2:0] = 3'b111;
      14'b01100101111100: pixel[2:0] = 3'b111;
      14'b01100101111101: pixel[2:0] = 3'b111;
      14'b01100101111110: pixel[2:0] = 3'b111;
      14'b01100101111111: pixel[2:0] = 3'b000;
      14'b01100110000000: pixel[2:0] = 3'b000;
      14'b01100110000001: pixel[2:0] = 3'b000;
      14'b01100110000010: pixel[2:0] = 3'b000;
      14'b01100110000011: pixel[2:0] = 3'b000;
      14'b01100110000100: pixel[2:0] = 3'b000;
      14'b01100110000101: pixel[2:0] = 3'b000;
      14'b01100110000110: pixel[2:0] = 3'b000;
      14'b01100110000111: pixel[2:0] = 3'b000;
      14'b01101000000000: pixel[2:0] = 3'b000;
      14'b01101000000001: pixel[2:0] = 3'b000;
      14'b01101000000010: pixel[2:0] = 3'b111;
      14'b01101000000011: pixel[2:0] = 3'b111;
      14'b01101000000100: pixel[2:0] = 3'b111;
      14'b01101000000101: pixel[2:0] = 3'b111;
      14'b01101000000110: pixel[2:0] = 3'b111;
      14'b01101000000111: pixel[2:0] = 3'b111;
      14'b01101000001000: pixel[2:0] = 3'b111;
      14'b01101000001001: pixel[2:0] = 3'b111;
      14'b01101000001010: pixel[2:0] = 3'b111;
      14'b01101000001011: pixel[2:0] = 3'b111;
      14'b01101000001100: pixel[2:0] = 3'b111;
      14'b01101000001101: pixel[2:0] = 3'b000;
      14'b01101000001110: pixel[2:0] = 3'b000;
      14'b01101000001111: pixel[2:0] = 3'b000;
      14'b01101000010000: pixel[2:0] = 3'b000;
      14'b01101000010001: pixel[2:0] = 3'b000;
      14'b01101000010010: pixel[2:0] = 3'b000;
      14'b01101000010011: pixel[2:0] = 3'b000;
      14'b01101000010100: pixel[2:0] = 3'b000;
      14'b01101000010101: pixel[2:0] = 3'b000;
      14'b01101000010110: pixel[2:0] = 3'b000;
      14'b01101000010111: pixel[2:0] = 3'b000;
      14'b01101000011000: pixel[2:0] = 3'b000;
      14'b01101000011001: pixel[2:0] = 3'b111;
      14'b01101000011010: pixel[2:0] = 3'b111;
      14'b01101000011011: pixel[2:0] = 3'b111;
      14'b01101000011100: pixel[2:0] = 3'b111;
      14'b01101000011101: pixel[2:0] = 3'b111;
      14'b01101000011110: pixel[2:0] = 3'b000;
      14'b01101000011111: pixel[2:0] = 3'b000;
      14'b01101000100000: pixel[2:0] = 3'b000;
      14'b01101000100001: pixel[2:0] = 3'b000;
      14'b01101000100010: pixel[2:0] = 3'b000;
      14'b01101000100011: pixel[2:0] = 3'b000;
      14'b01101000100100: pixel[2:0] = 3'b000;
      14'b01101000100101: pixel[2:0] = 3'b000;
      14'b01101000100110: pixel[2:0] = 3'b000;
      14'b01101000100111: pixel[2:0] = 3'b000;
      14'b01101000101000: pixel[2:0] = 3'b000;
      14'b01101000101001: pixel[2:0] = 3'b000;
      14'b01101000101010: pixel[2:0] = 3'b000;
      14'b01101000101011: pixel[2:0] = 3'b000;
      14'b01101000101100: pixel[2:0] = 3'b000;
      14'b01101000101101: pixel[2:0] = 3'b000;
      14'b01101000101110: pixel[2:0] = 3'b000;
      14'b01101000101111: pixel[2:0] = 3'b000;
      14'b01101000110000: pixel[2:0] = 3'b111;
      14'b01101000110001: pixel[2:0] = 3'b111;
      14'b01101000110010: pixel[2:0] = 3'b111;
      14'b01101000110011: pixel[2:0] = 3'b111;
      14'b01101000110100: pixel[2:0] = 3'b111;
      14'b01101000110101: pixel[2:0] = 3'b000;
      14'b01101000110110: pixel[2:0] = 3'b000;
      14'b01101000110111: pixel[2:0] = 3'b000;
      14'b01101000111000: pixel[2:0] = 3'b000;
      14'b01101000111001: pixel[2:0] = 3'b000;
      14'b01101000111010: pixel[2:0] = 3'b000;
      14'b01101000111011: pixel[2:0] = 3'b111;
      14'b01101000111100: pixel[2:0] = 3'b111;
      14'b01101000111101: pixel[2:0] = 3'b111;
      14'b01101000111110: pixel[2:0] = 3'b111;
      14'b01101000111111: pixel[2:0] = 3'b000;
      14'b01101001000000: pixel[2:0] = 3'b000;
      14'b01101001000001: pixel[2:0] = 3'b000;
      14'b01101001000010: pixel[2:0] = 3'b000;
      14'b01101001000011: pixel[2:0] = 3'b000;
      14'b01101001000100: pixel[2:0] = 3'b000;
      14'b01101001000101: pixel[2:0] = 3'b000;
      14'b01101001000110: pixel[2:0] = 3'b000;
      14'b01101001000111: pixel[2:0] = 3'b000;
      14'b01101001001000: pixel[2:0] = 3'b000;
      14'b01101001001001: pixel[2:0] = 3'b111;
      14'b01101001001010: pixel[2:0] = 3'b111;
      14'b01101001001011: pixel[2:0] = 3'b111;
      14'b01101001001100: pixel[2:0] = 3'b111;
      14'b01101001001101: pixel[2:0] = 3'b111;
      14'b01101001001110: pixel[2:0] = 3'b000;
      14'b01101001001111: pixel[2:0] = 3'b000;
      14'b01101001010000: pixel[2:0] = 3'b000;
      14'b01101001010001: pixel[2:0] = 3'b000;
      14'b01101001010010: pixel[2:0] = 3'b000;
      14'b01101001010011: pixel[2:0] = 3'b000;
      14'b01101001010100: pixel[2:0] = 3'b000;
      14'b01101001010101: pixel[2:0] = 3'b000;
      14'b01101001010110: pixel[2:0] = 3'b000;
      14'b01101001010111: pixel[2:0] = 3'b000;
      14'b01101001011000: pixel[2:0] = 3'b000;
      14'b01101001011001: pixel[2:0] = 3'b000;
      14'b01101001011010: pixel[2:0] = 3'b111;
      14'b01101001011011: pixel[2:0] = 3'b111;
      14'b01101001011100: pixel[2:0] = 3'b111;
      14'b01101001011101: pixel[2:0] = 3'b111;
      14'b01101001011110: pixel[2:0] = 3'b111;
      14'b01101001011111: pixel[2:0] = 3'b000;
      14'b01101001100000: pixel[2:0] = 3'b000;
      14'b01101001100001: pixel[2:0] = 3'b000;
      14'b01101001100010: pixel[2:0] = 3'b000;
      14'b01101001100011: pixel[2:0] = 3'b000;
      14'b01101001100100: pixel[2:0] = 3'b000;
      14'b01101001100101: pixel[2:0] = 3'b000;
      14'b01101001100110: pixel[2:0] = 3'b000;
      14'b01101001100111: pixel[2:0] = 3'b000;
      14'b01101001101000: pixel[2:0] = 3'b000;
      14'b01101001101001: pixel[2:0] = 3'b000;
      14'b01101001101010: pixel[2:0] = 3'b000;
      14'b01101001101011: pixel[2:0] = 3'b000;
      14'b01101001101100: pixel[2:0] = 3'b000;
      14'b01101001101101: pixel[2:0] = 3'b000;
      14'b01101001101110: pixel[2:0] = 3'b000;
      14'b01101001101111: pixel[2:0] = 3'b000;
      14'b01101001110000: pixel[2:0] = 3'b111;
      14'b01101001110001: pixel[2:0] = 3'b111;
      14'b01101001110010: pixel[2:0] = 3'b111;
      14'b01101001110011: pixel[2:0] = 3'b111;
      14'b01101001110100: pixel[2:0] = 3'b111;
      14'b01101001110101: pixel[2:0] = 3'b000;
      14'b01101001110110: pixel[2:0] = 3'b000;
      14'b01101001110111: pixel[2:0] = 3'b000;
      14'b01101001111000: pixel[2:0] = 3'b000;
      14'b01101001111001: pixel[2:0] = 3'b000;
      14'b01101001111010: pixel[2:0] = 3'b111;
      14'b01101001111011: pixel[2:0] = 3'b111;
      14'b01101001111100: pixel[2:0] = 3'b111;
      14'b01101001111101: pixel[2:0] = 3'b111;
      14'b01101001111110: pixel[2:0] = 3'b111;
      14'b01101001111111: pixel[2:0] = 3'b000;
      14'b01101010000000: pixel[2:0] = 3'b000;
      14'b01101010000001: pixel[2:0] = 3'b000;
      14'b01101010000010: pixel[2:0] = 3'b000;
      14'b01101010000011: pixel[2:0] = 3'b000;
      14'b01101010000100: pixel[2:0] = 3'b000;
      14'b01101010000101: pixel[2:0] = 3'b000;
      14'b01101010000110: pixel[2:0] = 3'b000;
      14'b01101010000111: pixel[2:0] = 3'b000;
      14'b01101100000000: pixel[2:0] = 3'b000;
      14'b01101100000001: pixel[2:0] = 3'b000;
      14'b01101100000010: pixel[2:0] = 3'b111;
      14'b01101100000011: pixel[2:0] = 3'b111;
      14'b01101100000100: pixel[2:0] = 3'b111;
      14'b01101100000101: pixel[2:0] = 3'b111;
      14'b01101100000110: pixel[2:0] = 3'b111;
      14'b01101100000111: pixel[2:0] = 3'b000;
      14'b01101100001000: pixel[2:0] = 3'b000;
      14'b01101100001001: pixel[2:0] = 3'b000;
      14'b01101100001010: pixel[2:0] = 3'b000;
      14'b01101100001011: pixel[2:0] = 3'b000;
      14'b01101100001100: pixel[2:0] = 3'b000;
      14'b01101100001101: pixel[2:0] = 3'b000;
      14'b01101100001110: pixel[2:0] = 3'b000;
      14'b01101100001111: pixel[2:0] = 3'b000;
      14'b01101100010000: pixel[2:0] = 3'b000;
      14'b01101100010001: pixel[2:0] = 3'b000;
      14'b01101100010010: pixel[2:0] = 3'b000;
      14'b01101100010011: pixel[2:0] = 3'b000;
      14'b01101100010100: pixel[2:0] = 3'b000;
      14'b01101100010101: pixel[2:0] = 3'b000;
      14'b01101100010110: pixel[2:0] = 3'b000;
      14'b01101100010111: pixel[2:0] = 3'b000;
      14'b01101100011000: pixel[2:0] = 3'b000;
      14'b01101100011001: pixel[2:0] = 3'b111;
      14'b01101100011010: pixel[2:0] = 3'b111;
      14'b01101100011011: pixel[2:0] = 3'b111;
      14'b01101100011100: pixel[2:0] = 3'b111;
      14'b01101100011101: pixel[2:0] = 3'b111;
      14'b01101100011110: pixel[2:0] = 3'b000;
      14'b01101100011111: pixel[2:0] = 3'b000;
      14'b01101100100000: pixel[2:0] = 3'b000;
      14'b01101100100001: pixel[2:0] = 3'b000;
      14'b01101100100010: pixel[2:0] = 3'b000;
      14'b01101100100011: pixel[2:0] = 3'b000;
      14'b01101100100100: pixel[2:0] = 3'b000;
      14'b01101100100101: pixel[2:0] = 3'b000;
      14'b01101100100110: pixel[2:0] = 3'b000;
      14'b01101100100111: pixel[2:0] = 3'b000;
      14'b01101100101000: pixel[2:0] = 3'b000;
      14'b01101100101001: pixel[2:0] = 3'b000;
      14'b01101100101010: pixel[2:0] = 3'b000;
      14'b01101100101011: pixel[2:0] = 3'b000;
      14'b01101100101100: pixel[2:0] = 3'b000;
      14'b01101100101101: pixel[2:0] = 3'b000;
      14'b01101100101110: pixel[2:0] = 3'b000;
      14'b01101100101111: pixel[2:0] = 3'b000;
      14'b01101100110000: pixel[2:0] = 3'b111;
      14'b01101100110001: pixel[2:0] = 3'b111;
      14'b01101100110010: pixel[2:0] = 3'b111;
      14'b01101100110011: pixel[2:0] = 3'b111;
      14'b01101100110100: pixel[2:0] = 3'b000;
      14'b01101100110101: pixel[2:0] = 3'b000;
      14'b01101100110110: pixel[2:0] = 3'b000;
      14'b01101100110111: pixel[2:0] = 3'b000;
      14'b01101100111000: pixel[2:0] = 3'b000;
      14'b01101100111001: pixel[2:0] = 3'b000;
      14'b01101100111010: pixel[2:0] = 3'b000;
      14'b01101100111011: pixel[2:0] = 3'b111;
      14'b01101100111100: pixel[2:0] = 3'b111;
      14'b01101100111101: pixel[2:0] = 3'b111;
      14'b01101100111110: pixel[2:0] = 3'b111;
      14'b01101100111111: pixel[2:0] = 3'b111;
      14'b01101101000000: pixel[2:0] = 3'b000;
      14'b01101101000001: pixel[2:0] = 3'b000;
      14'b01101101000010: pixel[2:0] = 3'b000;
      14'b01101101000011: pixel[2:0] = 3'b000;
      14'b01101101000100: pixel[2:0] = 3'b000;
      14'b01101101000101: pixel[2:0] = 3'b000;
      14'b01101101000110: pixel[2:0] = 3'b000;
      14'b01101101000111: pixel[2:0] = 3'b000;
      14'b01101101001000: pixel[2:0] = 3'b000;
      14'b01101101001001: pixel[2:0] = 3'b111;
      14'b01101101001010: pixel[2:0] = 3'b111;
      14'b01101101001011: pixel[2:0] = 3'b111;
      14'b01101101001100: pixel[2:0] = 3'b111;
      14'b01101101001101: pixel[2:0] = 3'b111;
      14'b01101101001110: pixel[2:0] = 3'b000;
      14'b01101101001111: pixel[2:0] = 3'b000;
      14'b01101101010000: pixel[2:0] = 3'b000;
      14'b01101101010001: pixel[2:0] = 3'b000;
      14'b01101101010010: pixel[2:0] = 3'b000;
      14'b01101101010011: pixel[2:0] = 3'b000;
      14'b01101101010100: pixel[2:0] = 3'b000;
      14'b01101101010101: pixel[2:0] = 3'b000;
      14'b01101101010110: pixel[2:0] = 3'b000;
      14'b01101101010111: pixel[2:0] = 3'b000;
      14'b01101101011000: pixel[2:0] = 3'b000;
      14'b01101101011001: pixel[2:0] = 3'b000;
      14'b01101101011010: pixel[2:0] = 3'b111;
      14'b01101101011011: pixel[2:0] = 3'b111;
      14'b01101101011100: pixel[2:0] = 3'b111;
      14'b01101101011101: pixel[2:0] = 3'b111;
      14'b01101101011110: pixel[2:0] = 3'b111;
      14'b01101101011111: pixel[2:0] = 3'b000;
      14'b01101101100000: pixel[2:0] = 3'b000;
      14'b01101101100001: pixel[2:0] = 3'b000;
      14'b01101101100010: pixel[2:0] = 3'b000;
      14'b01101101100011: pixel[2:0] = 3'b000;
      14'b01101101100100: pixel[2:0] = 3'b000;
      14'b01101101100101: pixel[2:0] = 3'b000;
      14'b01101101100110: pixel[2:0] = 3'b000;
      14'b01101101100111: pixel[2:0] = 3'b000;
      14'b01101101101000: pixel[2:0] = 3'b000;
      14'b01101101101001: pixel[2:0] = 3'b000;
      14'b01101101101010: pixel[2:0] = 3'b000;
      14'b01101101101011: pixel[2:0] = 3'b000;
      14'b01101101101100: pixel[2:0] = 3'b000;
      14'b01101101101101: pixel[2:0] = 3'b000;
      14'b01101101101110: pixel[2:0] = 3'b000;
      14'b01101101101111: pixel[2:0] = 3'b000;
      14'b01101101110000: pixel[2:0] = 3'b111;
      14'b01101101110001: pixel[2:0] = 3'b111;
      14'b01101101110010: pixel[2:0] = 3'b111;
      14'b01101101110011: pixel[2:0] = 3'b111;
      14'b01101101110100: pixel[2:0] = 3'b111;
      14'b01101101110101: pixel[2:0] = 3'b000;
      14'b01101101110110: pixel[2:0] = 3'b000;
      14'b01101101110111: pixel[2:0] = 3'b000;
      14'b01101101111000: pixel[2:0] = 3'b000;
      14'b01101101111001: pixel[2:0] = 3'b000;
      14'b01101101111010: pixel[2:0] = 3'b111;
      14'b01101101111011: pixel[2:0] = 3'b111;
      14'b01101101111100: pixel[2:0] = 3'b111;
      14'b01101101111101: pixel[2:0] = 3'b111;
      14'b01101101111110: pixel[2:0] = 3'b111;
      14'b01101101111111: pixel[2:0] = 3'b000;
      14'b01101110000000: pixel[2:0] = 3'b000;
      14'b01101110000001: pixel[2:0] = 3'b000;
      14'b01101110000010: pixel[2:0] = 3'b000;
      14'b01101110000011: pixel[2:0] = 3'b000;
      14'b01101110000100: pixel[2:0] = 3'b000;
      14'b01101110000101: pixel[2:0] = 3'b000;
      14'b01101110000110: pixel[2:0] = 3'b000;
      14'b01101110000111: pixel[2:0] = 3'b000;
      14'b01110000000000: pixel[2:0] = 3'b000;
      14'b01110000000001: pixel[2:0] = 3'b000;
      14'b01110000000010: pixel[2:0] = 3'b111;
      14'b01110000000011: pixel[2:0] = 3'b111;
      14'b01110000000100: pixel[2:0] = 3'b111;
      14'b01110000000101: pixel[2:0] = 3'b111;
      14'b01110000000110: pixel[2:0] = 3'b111;
      14'b01110000000111: pixel[2:0] = 3'b000;
      14'b01110000001000: pixel[2:0] = 3'b000;
      14'b01110000001001: pixel[2:0] = 3'b000;
      14'b01110000001010: pixel[2:0] = 3'b000;
      14'b01110000001011: pixel[2:0] = 3'b000;
      14'b01110000001100: pixel[2:0] = 3'b000;
      14'b01110000001101: pixel[2:0] = 3'b000;
      14'b01110000001110: pixel[2:0] = 3'b000;
      14'b01110000001111: pixel[2:0] = 3'b000;
      14'b01110000010000: pixel[2:0] = 3'b000;
      14'b01110000010001: pixel[2:0] = 3'b000;
      14'b01110000010010: pixel[2:0] = 3'b000;
      14'b01110000010011: pixel[2:0] = 3'b000;
      14'b01110000010100: pixel[2:0] = 3'b000;
      14'b01110000010101: pixel[2:0] = 3'b000;
      14'b01110000010110: pixel[2:0] = 3'b000;
      14'b01110000010111: pixel[2:0] = 3'b000;
      14'b01110000011000: pixel[2:0] = 3'b000;
      14'b01110000011001: pixel[2:0] = 3'b111;
      14'b01110000011010: pixel[2:0] = 3'b111;
      14'b01110000011011: pixel[2:0] = 3'b111;
      14'b01110000011100: pixel[2:0] = 3'b111;
      14'b01110000011101: pixel[2:0] = 3'b111;
      14'b01110000011110: pixel[2:0] = 3'b000;
      14'b01110000011111: pixel[2:0] = 3'b000;
      14'b01110000100000: pixel[2:0] = 3'b000;
      14'b01110000100001: pixel[2:0] = 3'b000;
      14'b01110000100010: pixel[2:0] = 3'b000;
      14'b01110000100011: pixel[2:0] = 3'b000;
      14'b01110000100100: pixel[2:0] = 3'b000;
      14'b01110000100101: pixel[2:0] = 3'b000;
      14'b01110000100110: pixel[2:0] = 3'b000;
      14'b01110000100111: pixel[2:0] = 3'b000;
      14'b01110000101000: pixel[2:0] = 3'b000;
      14'b01110000101001: pixel[2:0] = 3'b000;
      14'b01110000101010: pixel[2:0] = 3'b000;
      14'b01110000101011: pixel[2:0] = 3'b000;
      14'b01110000101100: pixel[2:0] = 3'b000;
      14'b01110000101101: pixel[2:0] = 3'b000;
      14'b01110000101110: pixel[2:0] = 3'b000;
      14'b01110000101111: pixel[2:0] = 3'b000;
      14'b01110000110000: pixel[2:0] = 3'b111;
      14'b01110000110001: pixel[2:0] = 3'b111;
      14'b01110000110010: pixel[2:0] = 3'b111;
      14'b01110000110011: pixel[2:0] = 3'b111;
      14'b01110000110100: pixel[2:0] = 3'b111;
      14'b01110000110101: pixel[2:0] = 3'b111;
      14'b01110000110110: pixel[2:0] = 3'b111;
      14'b01110000110111: pixel[2:0] = 3'b111;
      14'b01110000111000: pixel[2:0] = 3'b111;
      14'b01110000111001: pixel[2:0] = 3'b111;
      14'b01110000111010: pixel[2:0] = 3'b111;
      14'b01110000111011: pixel[2:0] = 3'b111;
      14'b01110000111100: pixel[2:0] = 3'b111;
      14'b01110000111101: pixel[2:0] = 3'b111;
      14'b01110000111110: pixel[2:0] = 3'b111;
      14'b01110000111111: pixel[2:0] = 3'b111;
      14'b01110001000000: pixel[2:0] = 3'b000;
      14'b01110001000001: pixel[2:0] = 3'b000;
      14'b01110001000010: pixel[2:0] = 3'b000;
      14'b01110001000011: pixel[2:0] = 3'b000;
      14'b01110001000100: pixel[2:0] = 3'b000;
      14'b01110001000101: pixel[2:0] = 3'b000;
      14'b01110001000110: pixel[2:0] = 3'b000;
      14'b01110001000111: pixel[2:0] = 3'b000;
      14'b01110001001000: pixel[2:0] = 3'b000;
      14'b01110001001001: pixel[2:0] = 3'b111;
      14'b01110001001010: pixel[2:0] = 3'b111;
      14'b01110001001011: pixel[2:0] = 3'b111;
      14'b01110001001100: pixel[2:0] = 3'b111;
      14'b01110001001101: pixel[2:0] = 3'b111;
      14'b01110001001110: pixel[2:0] = 3'b000;
      14'b01110001001111: pixel[2:0] = 3'b000;
      14'b01110001010000: pixel[2:0] = 3'b000;
      14'b01110001010001: pixel[2:0] = 3'b000;
      14'b01110001010010: pixel[2:0] = 3'b000;
      14'b01110001010011: pixel[2:0] = 3'b000;
      14'b01110001010100: pixel[2:0] = 3'b000;
      14'b01110001010101: pixel[2:0] = 3'b000;
      14'b01110001010110: pixel[2:0] = 3'b000;
      14'b01110001010111: pixel[2:0] = 3'b000;
      14'b01110001011000: pixel[2:0] = 3'b000;
      14'b01110001011001: pixel[2:0] = 3'b000;
      14'b01110001011010: pixel[2:0] = 3'b111;
      14'b01110001011011: pixel[2:0] = 3'b111;
      14'b01110001011100: pixel[2:0] = 3'b111;
      14'b01110001011101: pixel[2:0] = 3'b111;
      14'b01110001011110: pixel[2:0] = 3'b111;
      14'b01110001011111: pixel[2:0] = 3'b000;
      14'b01110001100000: pixel[2:0] = 3'b000;
      14'b01110001100001: pixel[2:0] = 3'b000;
      14'b01110001100010: pixel[2:0] = 3'b000;
      14'b01110001100011: pixel[2:0] = 3'b000;
      14'b01110001100100: pixel[2:0] = 3'b000;
      14'b01110001100101: pixel[2:0] = 3'b000;
      14'b01110001100110: pixel[2:0] = 3'b000;
      14'b01110001100111: pixel[2:0] = 3'b000;
      14'b01110001101000: pixel[2:0] = 3'b000;
      14'b01110001101001: pixel[2:0] = 3'b000;
      14'b01110001101010: pixel[2:0] = 3'b000;
      14'b01110001101011: pixel[2:0] = 3'b000;
      14'b01110001101100: pixel[2:0] = 3'b000;
      14'b01110001101101: pixel[2:0] = 3'b000;
      14'b01110001101110: pixel[2:0] = 3'b000;
      14'b01110001101111: pixel[2:0] = 3'b000;
      14'b01110001110000: pixel[2:0] = 3'b111;
      14'b01110001110001: pixel[2:0] = 3'b111;
      14'b01110001110010: pixel[2:0] = 3'b111;
      14'b01110001110011: pixel[2:0] = 3'b111;
      14'b01110001110100: pixel[2:0] = 3'b111;
      14'b01110001110101: pixel[2:0] = 3'b000;
      14'b01110001110110: pixel[2:0] = 3'b000;
      14'b01110001110111: pixel[2:0] = 3'b000;
      14'b01110001111000: pixel[2:0] = 3'b000;
      14'b01110001111001: pixel[2:0] = 3'b000;
      14'b01110001111010: pixel[2:0] = 3'b000;
      14'b01110001111011: pixel[2:0] = 3'b111;
      14'b01110001111100: pixel[2:0] = 3'b111;
      14'b01110001111101: pixel[2:0] = 3'b111;
      14'b01110001111110: pixel[2:0] = 3'b111;
      14'b01110001111111: pixel[2:0] = 3'b111;
      14'b01110010000000: pixel[2:0] = 3'b000;
      14'b01110010000001: pixel[2:0] = 3'b000;
      14'b01110010000010: pixel[2:0] = 3'b000;
      14'b01110010000011: pixel[2:0] = 3'b000;
      14'b01110010000100: pixel[2:0] = 3'b000;
      14'b01110010000101: pixel[2:0] = 3'b000;
      14'b01110010000110: pixel[2:0] = 3'b000;
      14'b01110010000111: pixel[2:0] = 3'b000;
      14'b01110100000000: pixel[2:0] = 3'b000;
      14'b01110100000001: pixel[2:0] = 3'b000;
      14'b01110100000010: pixel[2:0] = 3'b111;
      14'b01110100000011: pixel[2:0] = 3'b111;
      14'b01110100000100: pixel[2:0] = 3'b111;
      14'b01110100000101: pixel[2:0] = 3'b111;
      14'b01110100000110: pixel[2:0] = 3'b111;
      14'b01110100000111: pixel[2:0] = 3'b000;
      14'b01110100001000: pixel[2:0] = 3'b000;
      14'b01110100001001: pixel[2:0] = 3'b000;
      14'b01110100001010: pixel[2:0] = 3'b000;
      14'b01110100001011: pixel[2:0] = 3'b000;
      14'b01110100001100: pixel[2:0] = 3'b000;
      14'b01110100001101: pixel[2:0] = 3'b000;
      14'b01110100001110: pixel[2:0] = 3'b000;
      14'b01110100001111: pixel[2:0] = 3'b000;
      14'b01110100010000: pixel[2:0] = 3'b000;
      14'b01110100010001: pixel[2:0] = 3'b000;
      14'b01110100010010: pixel[2:0] = 3'b000;
      14'b01110100010011: pixel[2:0] = 3'b000;
      14'b01110100010100: pixel[2:0] = 3'b000;
      14'b01110100010101: pixel[2:0] = 3'b000;
      14'b01110100010110: pixel[2:0] = 3'b000;
      14'b01110100010111: pixel[2:0] = 3'b000;
      14'b01110100011000: pixel[2:0] = 3'b000;
      14'b01110100011001: pixel[2:0] = 3'b111;
      14'b01110100011010: pixel[2:0] = 3'b111;
      14'b01110100011011: pixel[2:0] = 3'b111;
      14'b01110100011100: pixel[2:0] = 3'b111;
      14'b01110100011101: pixel[2:0] = 3'b111;
      14'b01110100011110: pixel[2:0] = 3'b000;
      14'b01110100011111: pixel[2:0] = 3'b000;
      14'b01110100100000: pixel[2:0] = 3'b000;
      14'b01110100100001: pixel[2:0] = 3'b000;
      14'b01110100100010: pixel[2:0] = 3'b000;
      14'b01110100100011: pixel[2:0] = 3'b000;
      14'b01110100100100: pixel[2:0] = 3'b000;
      14'b01110100100101: pixel[2:0] = 3'b000;
      14'b01110100100110: pixel[2:0] = 3'b000;
      14'b01110100100111: pixel[2:0] = 3'b000;
      14'b01110100101000: pixel[2:0] = 3'b000;
      14'b01110100101001: pixel[2:0] = 3'b000;
      14'b01110100101010: pixel[2:0] = 3'b000;
      14'b01110100101011: pixel[2:0] = 3'b000;
      14'b01110100101100: pixel[2:0] = 3'b000;
      14'b01110100101101: pixel[2:0] = 3'b000;
      14'b01110100101110: pixel[2:0] = 3'b000;
      14'b01110100101111: pixel[2:0] = 3'b000;
      14'b01110100110000: pixel[2:0] = 3'b111;
      14'b01110100110001: pixel[2:0] = 3'b111;
      14'b01110100110010: pixel[2:0] = 3'b111;
      14'b01110100110011: pixel[2:0] = 3'b111;
      14'b01110100110100: pixel[2:0] = 3'b111;
      14'b01110100110101: pixel[2:0] = 3'b111;
      14'b01110100110110: pixel[2:0] = 3'b111;
      14'b01110100110111: pixel[2:0] = 3'b111;
      14'b01110100111000: pixel[2:0] = 3'b111;
      14'b01110100111001: pixel[2:0] = 3'b111;
      14'b01110100111010: pixel[2:0] = 3'b111;
      14'b01110100111011: pixel[2:0] = 3'b111;
      14'b01110100111100: pixel[2:0] = 3'b111;
      14'b01110100111101: pixel[2:0] = 3'b111;
      14'b01110100111110: pixel[2:0] = 3'b111;
      14'b01110100111111: pixel[2:0] = 3'b111;
      14'b01110101000000: pixel[2:0] = 3'b000;
      14'b01110101000001: pixel[2:0] = 3'b000;
      14'b01110101000010: pixel[2:0] = 3'b000;
      14'b01110101000011: pixel[2:0] = 3'b000;
      14'b01110101000100: pixel[2:0] = 3'b000;
      14'b01110101000101: pixel[2:0] = 3'b000;
      14'b01110101000110: pixel[2:0] = 3'b000;
      14'b01110101000111: pixel[2:0] = 3'b000;
      14'b01110101001000: pixel[2:0] = 3'b000;
      14'b01110101001001: pixel[2:0] = 3'b111;
      14'b01110101001010: pixel[2:0] = 3'b111;
      14'b01110101001011: pixel[2:0] = 3'b111;
      14'b01110101001100: pixel[2:0] = 3'b111;
      14'b01110101001101: pixel[2:0] = 3'b111;
      14'b01110101001110: pixel[2:0] = 3'b000;
      14'b01110101001111: pixel[2:0] = 3'b000;
      14'b01110101010000: pixel[2:0] = 3'b000;
      14'b01110101010001: pixel[2:0] = 3'b000;
      14'b01110101010010: pixel[2:0] = 3'b000;
      14'b01110101010011: pixel[2:0] = 3'b000;
      14'b01110101010100: pixel[2:0] = 3'b000;
      14'b01110101010101: pixel[2:0] = 3'b000;
      14'b01110101010110: pixel[2:0] = 3'b000;
      14'b01110101010111: pixel[2:0] = 3'b000;
      14'b01110101011000: pixel[2:0] = 3'b000;
      14'b01110101011001: pixel[2:0] = 3'b000;
      14'b01110101011010: pixel[2:0] = 3'b111;
      14'b01110101011011: pixel[2:0] = 3'b111;
      14'b01110101011100: pixel[2:0] = 3'b111;
      14'b01110101011101: pixel[2:0] = 3'b111;
      14'b01110101011110: pixel[2:0] = 3'b111;
      14'b01110101011111: pixel[2:0] = 3'b000;
      14'b01110101100000: pixel[2:0] = 3'b000;
      14'b01110101100001: pixel[2:0] = 3'b000;
      14'b01110101100010: pixel[2:0] = 3'b000;
      14'b01110101100011: pixel[2:0] = 3'b000;
      14'b01110101100100: pixel[2:0] = 3'b000;
      14'b01110101100101: pixel[2:0] = 3'b000;
      14'b01110101100110: pixel[2:0] = 3'b000;
      14'b01110101100111: pixel[2:0] = 3'b000;
      14'b01110101101000: pixel[2:0] = 3'b000;
      14'b01110101101001: pixel[2:0] = 3'b000;
      14'b01110101101010: pixel[2:0] = 3'b000;
      14'b01110101101011: pixel[2:0] = 3'b000;
      14'b01110101101100: pixel[2:0] = 3'b000;
      14'b01110101101101: pixel[2:0] = 3'b000;
      14'b01110101101110: pixel[2:0] = 3'b000;
      14'b01110101101111: pixel[2:0] = 3'b000;
      14'b01110101110000: pixel[2:0] = 3'b111;
      14'b01110101110001: pixel[2:0] = 3'b111;
      14'b01110101110010: pixel[2:0] = 3'b111;
      14'b01110101110011: pixel[2:0] = 3'b111;
      14'b01110101110100: pixel[2:0] = 3'b111;
      14'b01110101110101: pixel[2:0] = 3'b000;
      14'b01110101110110: pixel[2:0] = 3'b000;
      14'b01110101110111: pixel[2:0] = 3'b000;
      14'b01110101111000: pixel[2:0] = 3'b000;
      14'b01110101111001: pixel[2:0] = 3'b000;
      14'b01110101111010: pixel[2:0] = 3'b000;
      14'b01110101111011: pixel[2:0] = 3'b111;
      14'b01110101111100: pixel[2:0] = 3'b111;
      14'b01110101111101: pixel[2:0] = 3'b111;
      14'b01110101111110: pixel[2:0] = 3'b111;
      14'b01110101111111: pixel[2:0] = 3'b111;
      14'b01110110000000: pixel[2:0] = 3'b000;
      14'b01110110000001: pixel[2:0] = 3'b000;
      14'b01110110000010: pixel[2:0] = 3'b000;
      14'b01110110000011: pixel[2:0] = 3'b000;
      14'b01110110000100: pixel[2:0] = 3'b000;
      14'b01110110000101: pixel[2:0] = 3'b000;
      14'b01110110000110: pixel[2:0] = 3'b000;
      14'b01110110000111: pixel[2:0] = 3'b000;
      14'b01111000000000: pixel[2:0] = 3'b000;
      14'b01111000000001: pixel[2:0] = 3'b000;
      14'b01111000000010: pixel[2:0] = 3'b111;
      14'b01111000000011: pixel[2:0] = 3'b111;
      14'b01111000000100: pixel[2:0] = 3'b111;
      14'b01111000000101: pixel[2:0] = 3'b111;
      14'b01111000000110: pixel[2:0] = 3'b111;
      14'b01111000000111: pixel[2:0] = 3'b000;
      14'b01111000001000: pixel[2:0] = 3'b000;
      14'b01111000001001: pixel[2:0] = 3'b000;
      14'b01111000001010: pixel[2:0] = 3'b000;
      14'b01111000001011: pixel[2:0] = 3'b000;
      14'b01111000001100: pixel[2:0] = 3'b000;
      14'b01111000001101: pixel[2:0] = 3'b000;
      14'b01111000001110: pixel[2:0] = 3'b000;
      14'b01111000001111: pixel[2:0] = 3'b000;
      14'b01111000010000: pixel[2:0] = 3'b000;
      14'b01111000010001: pixel[2:0] = 3'b000;
      14'b01111000010010: pixel[2:0] = 3'b000;
      14'b01111000010011: pixel[2:0] = 3'b000;
      14'b01111000010100: pixel[2:0] = 3'b000;
      14'b01111000010101: pixel[2:0] = 3'b000;
      14'b01111000010110: pixel[2:0] = 3'b000;
      14'b01111000010111: pixel[2:0] = 3'b000;
      14'b01111000011000: pixel[2:0] = 3'b000;
      14'b01111000011001: pixel[2:0] = 3'b111;
      14'b01111000011010: pixel[2:0] = 3'b111;
      14'b01111000011011: pixel[2:0] = 3'b111;
      14'b01111000011100: pixel[2:0] = 3'b111;
      14'b01111000011101: pixel[2:0] = 3'b111;
      14'b01111000011110: pixel[2:0] = 3'b000;
      14'b01111000011111: pixel[2:0] = 3'b000;
      14'b01111000100000: pixel[2:0] = 3'b000;
      14'b01111000100001: pixel[2:0] = 3'b000;
      14'b01111000100010: pixel[2:0] = 3'b000;
      14'b01111000100011: pixel[2:0] = 3'b000;
      14'b01111000100100: pixel[2:0] = 3'b000;
      14'b01111000100101: pixel[2:0] = 3'b000;
      14'b01111000100110: pixel[2:0] = 3'b000;
      14'b01111000100111: pixel[2:0] = 3'b000;
      14'b01111000101000: pixel[2:0] = 3'b000;
      14'b01111000101001: pixel[2:0] = 3'b000;
      14'b01111000101010: pixel[2:0] = 3'b000;
      14'b01111000101011: pixel[2:0] = 3'b000;
      14'b01111000101100: pixel[2:0] = 3'b000;
      14'b01111000101101: pixel[2:0] = 3'b000;
      14'b01111000101110: pixel[2:0] = 3'b000;
      14'b01111000101111: pixel[2:0] = 3'b111;
      14'b01111000110000: pixel[2:0] = 3'b111;
      14'b01111000110001: pixel[2:0] = 3'b111;
      14'b01111000110010: pixel[2:0] = 3'b111;
      14'b01111000110011: pixel[2:0] = 3'b111;
      14'b01111000110100: pixel[2:0] = 3'b111;
      14'b01111000110101: pixel[2:0] = 3'b111;
      14'b01111000110110: pixel[2:0] = 3'b111;
      14'b01111000110111: pixel[2:0] = 3'b111;
      14'b01111000111000: pixel[2:0] = 3'b111;
      14'b01111000111001: pixel[2:0] = 3'b111;
      14'b01111000111010: pixel[2:0] = 3'b111;
      14'b01111000111011: pixel[2:0] = 3'b111;
      14'b01111000111100: pixel[2:0] = 3'b111;
      14'b01111000111101: pixel[2:0] = 3'b111;
      14'b01111000111110: pixel[2:0] = 3'b111;
      14'b01111000111111: pixel[2:0] = 3'b111;
      14'b01111001000000: pixel[2:0] = 3'b000;
      14'b01111001000001: pixel[2:0] = 3'b000;
      14'b01111001000010: pixel[2:0] = 3'b000;
      14'b01111001000011: pixel[2:0] = 3'b000;
      14'b01111001000100: pixel[2:0] = 3'b000;
      14'b01111001000101: pixel[2:0] = 3'b000;
      14'b01111001000110: pixel[2:0] = 3'b000;
      14'b01111001000111: pixel[2:0] = 3'b000;
      14'b01111001001000: pixel[2:0] = 3'b000;
      14'b01111001001001: pixel[2:0] = 3'b111;
      14'b01111001001010: pixel[2:0] = 3'b111;
      14'b01111001001011: pixel[2:0] = 3'b111;
      14'b01111001001100: pixel[2:0] = 3'b111;
      14'b01111001001101: pixel[2:0] = 3'b111;
      14'b01111001001110: pixel[2:0] = 3'b000;
      14'b01111001001111: pixel[2:0] = 3'b000;
      14'b01111001010000: pixel[2:0] = 3'b000;
      14'b01111001010001: pixel[2:0] = 3'b000;
      14'b01111001010010: pixel[2:0] = 3'b000;
      14'b01111001010011: pixel[2:0] = 3'b000;
      14'b01111001010100: pixel[2:0] = 3'b000;
      14'b01111001010101: pixel[2:0] = 3'b000;
      14'b01111001010110: pixel[2:0] = 3'b000;
      14'b01111001010111: pixel[2:0] = 3'b000;
      14'b01111001011000: pixel[2:0] = 3'b000;
      14'b01111001011001: pixel[2:0] = 3'b000;
      14'b01111001011010: pixel[2:0] = 3'b111;
      14'b01111001011011: pixel[2:0] = 3'b111;
      14'b01111001011100: pixel[2:0] = 3'b111;
      14'b01111001011101: pixel[2:0] = 3'b111;
      14'b01111001011110: pixel[2:0] = 3'b111;
      14'b01111001011111: pixel[2:0] = 3'b000;
      14'b01111001100000: pixel[2:0] = 3'b000;
      14'b01111001100001: pixel[2:0] = 3'b000;
      14'b01111001100010: pixel[2:0] = 3'b000;
      14'b01111001100011: pixel[2:0] = 3'b000;
      14'b01111001100100: pixel[2:0] = 3'b000;
      14'b01111001100101: pixel[2:0] = 3'b000;
      14'b01111001100110: pixel[2:0] = 3'b000;
      14'b01111001100111: pixel[2:0] = 3'b000;
      14'b01111001101000: pixel[2:0] = 3'b000;
      14'b01111001101001: pixel[2:0] = 3'b000;
      14'b01111001101010: pixel[2:0] = 3'b000;
      14'b01111001101011: pixel[2:0] = 3'b000;
      14'b01111001101100: pixel[2:0] = 3'b000;
      14'b01111001101101: pixel[2:0] = 3'b000;
      14'b01111001101110: pixel[2:0] = 3'b000;
      14'b01111001101111: pixel[2:0] = 3'b000;
      14'b01111001110000: pixel[2:0] = 3'b111;
      14'b01111001110001: pixel[2:0] = 3'b111;
      14'b01111001110010: pixel[2:0] = 3'b111;
      14'b01111001110011: pixel[2:0] = 3'b111;
      14'b01111001110100: pixel[2:0] = 3'b111;
      14'b01111001110101: pixel[2:0] = 3'b000;
      14'b01111001110110: pixel[2:0] = 3'b000;
      14'b01111001110111: pixel[2:0] = 3'b000;
      14'b01111001111000: pixel[2:0] = 3'b000;
      14'b01111001111001: pixel[2:0] = 3'b000;
      14'b01111001111010: pixel[2:0] = 3'b000;
      14'b01111001111011: pixel[2:0] = 3'b111;
      14'b01111001111100: pixel[2:0] = 3'b111;
      14'b01111001111101: pixel[2:0] = 3'b111;
      14'b01111001111110: pixel[2:0] = 3'b111;
      14'b01111001111111: pixel[2:0] = 3'b111;
      14'b01111010000000: pixel[2:0] = 3'b000;
      14'b01111010000001: pixel[2:0] = 3'b000;
      14'b01111010000010: pixel[2:0] = 3'b000;
      14'b01111010000011: pixel[2:0] = 3'b000;
      14'b01111010000100: pixel[2:0] = 3'b000;
      14'b01111010000101: pixel[2:0] = 3'b000;
      14'b01111010000110: pixel[2:0] = 3'b000;
      14'b01111010000111: pixel[2:0] = 3'b000;
      14'b01111100000000: pixel[2:0] = 3'b000;
      14'b01111100000001: pixel[2:0] = 3'b000;
      14'b01111100000010: pixel[2:0] = 3'b111;
      14'b01111100000011: pixel[2:0] = 3'b111;
      14'b01111100000100: pixel[2:0] = 3'b111;
      14'b01111100000101: pixel[2:0] = 3'b111;
      14'b01111100000110: pixel[2:0] = 3'b111;
      14'b01111100000111: pixel[2:0] = 3'b000;
      14'b01111100001000: pixel[2:0] = 3'b000;
      14'b01111100001001: pixel[2:0] = 3'b000;
      14'b01111100001010: pixel[2:0] = 3'b000;
      14'b01111100001011: pixel[2:0] = 3'b000;
      14'b01111100001100: pixel[2:0] = 3'b000;
      14'b01111100001101: pixel[2:0] = 3'b000;
      14'b01111100001110: pixel[2:0] = 3'b000;
      14'b01111100001111: pixel[2:0] = 3'b000;
      14'b01111100010000: pixel[2:0] = 3'b000;
      14'b01111100010001: pixel[2:0] = 3'b000;
      14'b01111100010010: pixel[2:0] = 3'b000;
      14'b01111100010011: pixel[2:0] = 3'b000;
      14'b01111100010100: pixel[2:0] = 3'b000;
      14'b01111100010101: pixel[2:0] = 3'b000;
      14'b01111100010110: pixel[2:0] = 3'b000;
      14'b01111100010111: pixel[2:0] = 3'b000;
      14'b01111100011000: pixel[2:0] = 3'b000;
      14'b01111100011001: pixel[2:0] = 3'b111;
      14'b01111100011010: pixel[2:0] = 3'b111;
      14'b01111100011011: pixel[2:0] = 3'b111;
      14'b01111100011100: pixel[2:0] = 3'b111;
      14'b01111100011101: pixel[2:0] = 3'b111;
      14'b01111100011110: pixel[2:0] = 3'b000;
      14'b01111100011111: pixel[2:0] = 3'b000;
      14'b01111100100000: pixel[2:0] = 3'b000;
      14'b01111100100001: pixel[2:0] = 3'b000;
      14'b01111100100010: pixel[2:0] = 3'b000;
      14'b01111100100011: pixel[2:0] = 3'b000;
      14'b01111100100100: pixel[2:0] = 3'b000;
      14'b01111100100101: pixel[2:0] = 3'b000;
      14'b01111100100110: pixel[2:0] = 3'b000;
      14'b01111100100111: pixel[2:0] = 3'b000;
      14'b01111100101000: pixel[2:0] = 3'b000;
      14'b01111100101001: pixel[2:0] = 3'b000;
      14'b01111100101010: pixel[2:0] = 3'b000;
      14'b01111100101011: pixel[2:0] = 3'b000;
      14'b01111100101100: pixel[2:0] = 3'b000;
      14'b01111100101101: pixel[2:0] = 3'b000;
      14'b01111100101110: pixel[2:0] = 3'b000;
      14'b01111100101111: pixel[2:0] = 3'b111;
      14'b01111100110000: pixel[2:0] = 3'b111;
      14'b01111100110001: pixel[2:0] = 3'b111;
      14'b01111100110010: pixel[2:0] = 3'b111;
      14'b01111100110011: pixel[2:0] = 3'b111;
      14'b01111100110100: pixel[2:0] = 3'b111;
      14'b01111100110101: pixel[2:0] = 3'b111;
      14'b01111100110110: pixel[2:0] = 3'b111;
      14'b01111100110111: pixel[2:0] = 3'b111;
      14'b01111100111000: pixel[2:0] = 3'b111;
      14'b01111100111001: pixel[2:0] = 3'b111;
      14'b01111100111010: pixel[2:0] = 3'b111;
      14'b01111100111011: pixel[2:0] = 3'b111;
      14'b01111100111100: pixel[2:0] = 3'b111;
      14'b01111100111101: pixel[2:0] = 3'b111;
      14'b01111100111110: pixel[2:0] = 3'b111;
      14'b01111100111111: pixel[2:0] = 3'b111;
      14'b01111101000000: pixel[2:0] = 3'b000;
      14'b01111101000001: pixel[2:0] = 3'b000;
      14'b01111101000010: pixel[2:0] = 3'b000;
      14'b01111101000011: pixel[2:0] = 3'b000;
      14'b01111101000100: pixel[2:0] = 3'b000;
      14'b01111101000101: pixel[2:0] = 3'b000;
      14'b01111101000110: pixel[2:0] = 3'b000;
      14'b01111101000111: pixel[2:0] = 3'b000;
      14'b01111101001000: pixel[2:0] = 3'b000;
      14'b01111101001001: pixel[2:0] = 3'b111;
      14'b01111101001010: pixel[2:0] = 3'b111;
      14'b01111101001011: pixel[2:0] = 3'b111;
      14'b01111101001100: pixel[2:0] = 3'b111;
      14'b01111101001101: pixel[2:0] = 3'b111;
      14'b01111101001110: pixel[2:0] = 3'b000;
      14'b01111101001111: pixel[2:0] = 3'b000;
      14'b01111101010000: pixel[2:0] = 3'b000;
      14'b01111101010001: pixel[2:0] = 3'b000;
      14'b01111101010010: pixel[2:0] = 3'b000;
      14'b01111101010011: pixel[2:0] = 3'b000;
      14'b01111101010100: pixel[2:0] = 3'b000;
      14'b01111101010101: pixel[2:0] = 3'b000;
      14'b01111101010110: pixel[2:0] = 3'b000;
      14'b01111101010111: pixel[2:0] = 3'b000;
      14'b01111101011000: pixel[2:0] = 3'b000;
      14'b01111101011001: pixel[2:0] = 3'b000;
      14'b01111101011010: pixel[2:0] = 3'b111;
      14'b01111101011011: pixel[2:0] = 3'b111;
      14'b01111101011100: pixel[2:0] = 3'b111;
      14'b01111101011101: pixel[2:0] = 3'b111;
      14'b01111101011110: pixel[2:0] = 3'b111;
      14'b01111101011111: pixel[2:0] = 3'b000;
      14'b01111101100000: pixel[2:0] = 3'b000;
      14'b01111101100001: pixel[2:0] = 3'b000;
      14'b01111101100010: pixel[2:0] = 3'b000;
      14'b01111101100011: pixel[2:0] = 3'b000;
      14'b01111101100100: pixel[2:0] = 3'b000;
      14'b01111101100101: pixel[2:0] = 3'b000;
      14'b01111101100110: pixel[2:0] = 3'b000;
      14'b01111101100111: pixel[2:0] = 3'b000;
      14'b01111101101000: pixel[2:0] = 3'b000;
      14'b01111101101001: pixel[2:0] = 3'b000;
      14'b01111101101010: pixel[2:0] = 3'b000;
      14'b01111101101011: pixel[2:0] = 3'b000;
      14'b01111101101100: pixel[2:0] = 3'b000;
      14'b01111101101101: pixel[2:0] = 3'b000;
      14'b01111101101110: pixel[2:0] = 3'b000;
      14'b01111101101111: pixel[2:0] = 3'b000;
      14'b01111101110000: pixel[2:0] = 3'b111;
      14'b01111101110001: pixel[2:0] = 3'b111;
      14'b01111101110010: pixel[2:0] = 3'b111;
      14'b01111101110011: pixel[2:0] = 3'b111;
      14'b01111101110100: pixel[2:0] = 3'b111;
      14'b01111101110101: pixel[2:0] = 3'b000;
      14'b01111101110110: pixel[2:0] = 3'b000;
      14'b01111101110111: pixel[2:0] = 3'b000;
      14'b01111101111000: pixel[2:0] = 3'b000;
      14'b01111101111001: pixel[2:0] = 3'b000;
      14'b01111101111010: pixel[2:0] = 3'b000;
      14'b01111101111011: pixel[2:0] = 3'b000;
      14'b01111101111100: pixel[2:0] = 3'b111;
      14'b01111101111101: pixel[2:0] = 3'b111;
      14'b01111101111110: pixel[2:0] = 3'b111;
      14'b01111101111111: pixel[2:0] = 3'b111;
      14'b01111110000000: pixel[2:0] = 3'b111;
      14'b01111110000001: pixel[2:0] = 3'b000;
      14'b01111110000010: pixel[2:0] = 3'b000;
      14'b01111110000011: pixel[2:0] = 3'b000;
      14'b01111110000100: pixel[2:0] = 3'b000;
      14'b01111110000101: pixel[2:0] = 3'b000;
      14'b01111110000110: pixel[2:0] = 3'b000;
      14'b01111110000111: pixel[2:0] = 3'b000;
      14'b10000000000000: pixel[2:0] = 3'b000;
      14'b10000000000001: pixel[2:0] = 3'b000;
      14'b10000000000010: pixel[2:0] = 3'b111;
      14'b10000000000011: pixel[2:0] = 3'b111;
      14'b10000000000100: pixel[2:0] = 3'b111;
      14'b10000000000101: pixel[2:0] = 3'b111;
      14'b10000000000110: pixel[2:0] = 3'b111;
      14'b10000000000111: pixel[2:0] = 3'b000;
      14'b10000000001000: pixel[2:0] = 3'b000;
      14'b10000000001001: pixel[2:0] = 3'b000;
      14'b10000000001010: pixel[2:0] = 3'b000;
      14'b10000000001011: pixel[2:0] = 3'b000;
      14'b10000000001100: pixel[2:0] = 3'b000;
      14'b10000000001101: pixel[2:0] = 3'b000;
      14'b10000000001110: pixel[2:0] = 3'b000;
      14'b10000000001111: pixel[2:0] = 3'b000;
      14'b10000000010000: pixel[2:0] = 3'b000;
      14'b10000000010001: pixel[2:0] = 3'b000;
      14'b10000000010010: pixel[2:0] = 3'b000;
      14'b10000000010011: pixel[2:0] = 3'b000;
      14'b10000000010100: pixel[2:0] = 3'b000;
      14'b10000000010101: pixel[2:0] = 3'b000;
      14'b10000000010110: pixel[2:0] = 3'b000;
      14'b10000000010111: pixel[2:0] = 3'b000;
      14'b10000000011000: pixel[2:0] = 3'b000;
      14'b10000000011001: pixel[2:0] = 3'b111;
      14'b10000000011010: pixel[2:0] = 3'b111;
      14'b10000000011011: pixel[2:0] = 3'b111;
      14'b10000000011100: pixel[2:0] = 3'b111;
      14'b10000000011101: pixel[2:0] = 3'b111;
      14'b10000000011110: pixel[2:0] = 3'b000;
      14'b10000000011111: pixel[2:0] = 3'b000;
      14'b10000000100000: pixel[2:0] = 3'b000;
      14'b10000000100001: pixel[2:0] = 3'b000;
      14'b10000000100010: pixel[2:0] = 3'b000;
      14'b10000000100011: pixel[2:0] = 3'b000;
      14'b10000000100100: pixel[2:0] = 3'b000;
      14'b10000000100101: pixel[2:0] = 3'b000;
      14'b10000000100110: pixel[2:0] = 3'b000;
      14'b10000000100111: pixel[2:0] = 3'b000;
      14'b10000000101000: pixel[2:0] = 3'b000;
      14'b10000000101001: pixel[2:0] = 3'b000;
      14'b10000000101010: pixel[2:0] = 3'b000;
      14'b10000000101011: pixel[2:0] = 3'b000;
      14'b10000000101100: pixel[2:0] = 3'b000;
      14'b10000000101101: pixel[2:0] = 3'b000;
      14'b10000000101110: pixel[2:0] = 3'b000;
      14'b10000000101111: pixel[2:0] = 3'b111;
      14'b10000000110000: pixel[2:0] = 3'b111;
      14'b10000000110001: pixel[2:0] = 3'b111;
      14'b10000000110010: pixel[2:0] = 3'b111;
      14'b10000000110011: pixel[2:0] = 3'b111;
      14'b10000000110100: pixel[2:0] = 3'b111;
      14'b10000000110101: pixel[2:0] = 3'b111;
      14'b10000000110110: pixel[2:0] = 3'b111;
      14'b10000000110111: pixel[2:0] = 3'b111;
      14'b10000000111000: pixel[2:0] = 3'b111;
      14'b10000000111001: pixel[2:0] = 3'b111;
      14'b10000000111010: pixel[2:0] = 3'b111;
      14'b10000000111011: pixel[2:0] = 3'b111;
      14'b10000000111100: pixel[2:0] = 3'b111;
      14'b10000000111101: pixel[2:0] = 3'b111;
      14'b10000000111110: pixel[2:0] = 3'b111;
      14'b10000000111111: pixel[2:0] = 3'b111;
      14'b10000001000000: pixel[2:0] = 3'b111;
      14'b10000001000001: pixel[2:0] = 3'b000;
      14'b10000001000010: pixel[2:0] = 3'b000;
      14'b10000001000011: pixel[2:0] = 3'b000;
      14'b10000001000100: pixel[2:0] = 3'b000;
      14'b10000001000101: pixel[2:0] = 3'b000;
      14'b10000001000110: pixel[2:0] = 3'b000;
      14'b10000001000111: pixel[2:0] = 3'b000;
      14'b10000001001000: pixel[2:0] = 3'b000;
      14'b10000001001001: pixel[2:0] = 3'b111;
      14'b10000001001010: pixel[2:0] = 3'b111;
      14'b10000001001011: pixel[2:0] = 3'b111;
      14'b10000001001100: pixel[2:0] = 3'b111;
      14'b10000001001101: pixel[2:0] = 3'b111;
      14'b10000001001110: pixel[2:0] = 3'b000;
      14'b10000001001111: pixel[2:0] = 3'b000;
      14'b10000001010000: pixel[2:0] = 3'b000;
      14'b10000001010001: pixel[2:0] = 3'b000;
      14'b10000001010010: pixel[2:0] = 3'b000;
      14'b10000001010011: pixel[2:0] = 3'b000;
      14'b10000001010100: pixel[2:0] = 3'b000;
      14'b10000001010101: pixel[2:0] = 3'b000;
      14'b10000001010110: pixel[2:0] = 3'b000;
      14'b10000001010111: pixel[2:0] = 3'b000;
      14'b10000001011000: pixel[2:0] = 3'b000;
      14'b10000001011001: pixel[2:0] = 3'b000;
      14'b10000001011010: pixel[2:0] = 3'b111;
      14'b10000001011011: pixel[2:0] = 3'b111;
      14'b10000001011100: pixel[2:0] = 3'b111;
      14'b10000001011101: pixel[2:0] = 3'b111;
      14'b10000001011110: pixel[2:0] = 3'b111;
      14'b10000001011111: pixel[2:0] = 3'b000;
      14'b10000001100000: pixel[2:0] = 3'b000;
      14'b10000001100001: pixel[2:0] = 3'b000;
      14'b10000001100010: pixel[2:0] = 3'b000;
      14'b10000001100011: pixel[2:0] = 3'b000;
      14'b10000001100100: pixel[2:0] = 3'b000;
      14'b10000001100101: pixel[2:0] = 3'b000;
      14'b10000001100110: pixel[2:0] = 3'b000;
      14'b10000001100111: pixel[2:0] = 3'b000;
      14'b10000001101000: pixel[2:0] = 3'b000;
      14'b10000001101001: pixel[2:0] = 3'b000;
      14'b10000001101010: pixel[2:0] = 3'b000;
      14'b10000001101011: pixel[2:0] = 3'b000;
      14'b10000001101100: pixel[2:0] = 3'b000;
      14'b10000001101101: pixel[2:0] = 3'b000;
      14'b10000001101110: pixel[2:0] = 3'b000;
      14'b10000001101111: pixel[2:0] = 3'b000;
      14'b10000001110000: pixel[2:0] = 3'b111;
      14'b10000001110001: pixel[2:0] = 3'b111;
      14'b10000001110010: pixel[2:0] = 3'b111;
      14'b10000001110011: pixel[2:0] = 3'b111;
      14'b10000001110100: pixel[2:0] = 3'b111;
      14'b10000001110101: pixel[2:0] = 3'b000;
      14'b10000001110110: pixel[2:0] = 3'b000;
      14'b10000001110111: pixel[2:0] = 3'b000;
      14'b10000001111000: pixel[2:0] = 3'b000;
      14'b10000001111001: pixel[2:0] = 3'b000;
      14'b10000001111010: pixel[2:0] = 3'b000;
      14'b10000001111011: pixel[2:0] = 3'b000;
      14'b10000001111100: pixel[2:0] = 3'b111;
      14'b10000001111101: pixel[2:0] = 3'b111;
      14'b10000001111110: pixel[2:0] = 3'b111;
      14'b10000001111111: pixel[2:0] = 3'b111;
      14'b10000010000000: pixel[2:0] = 3'b111;
      14'b10000010000001: pixel[2:0] = 3'b000;
      14'b10000010000010: pixel[2:0] = 3'b000;
      14'b10000010000011: pixel[2:0] = 3'b000;
      14'b10000010000100: pixel[2:0] = 3'b000;
      14'b10000010000101: pixel[2:0] = 3'b000;
      14'b10000010000110: pixel[2:0] = 3'b000;
      14'b10000010000111: pixel[2:0] = 3'b000;
      14'b10000100000000: pixel[2:0] = 3'b000;
      14'b10000100000001: pixel[2:0] = 3'b000;
      14'b10000100000010: pixel[2:0] = 3'b111;
      14'b10000100000011: pixel[2:0] = 3'b111;
      14'b10000100000100: pixel[2:0] = 3'b111;
      14'b10000100000101: pixel[2:0] = 3'b111;
      14'b10000100000110: pixel[2:0] = 3'b111;
      14'b10000100000111: pixel[2:0] = 3'b000;
      14'b10000100001000: pixel[2:0] = 3'b000;
      14'b10000100001001: pixel[2:0] = 3'b000;
      14'b10000100001010: pixel[2:0] = 3'b000;
      14'b10000100001011: pixel[2:0] = 3'b000;
      14'b10000100001100: pixel[2:0] = 3'b000;
      14'b10000100001101: pixel[2:0] = 3'b000;
      14'b10000100001110: pixel[2:0] = 3'b000;
      14'b10000100001111: pixel[2:0] = 3'b000;
      14'b10000100010000: pixel[2:0] = 3'b000;
      14'b10000100010001: pixel[2:0] = 3'b000;
      14'b10000100010010: pixel[2:0] = 3'b000;
      14'b10000100010011: pixel[2:0] = 3'b000;
      14'b10000100010100: pixel[2:0] = 3'b000;
      14'b10000100010101: pixel[2:0] = 3'b000;
      14'b10000100010110: pixel[2:0] = 3'b000;
      14'b10000100010111: pixel[2:0] = 3'b000;
      14'b10000100011000: pixel[2:0] = 3'b000;
      14'b10000100011001: pixel[2:0] = 3'b111;
      14'b10000100011010: pixel[2:0] = 3'b111;
      14'b10000100011011: pixel[2:0] = 3'b111;
      14'b10000100011100: pixel[2:0] = 3'b111;
      14'b10000100011101: pixel[2:0] = 3'b111;
      14'b10000100011110: pixel[2:0] = 3'b000;
      14'b10000100011111: pixel[2:0] = 3'b000;
      14'b10000100100000: pixel[2:0] = 3'b000;
      14'b10000100100001: pixel[2:0] = 3'b000;
      14'b10000100100010: pixel[2:0] = 3'b000;
      14'b10000100100011: pixel[2:0] = 3'b000;
      14'b10000100100100: pixel[2:0] = 3'b000;
      14'b10000100100101: pixel[2:0] = 3'b000;
      14'b10000100100110: pixel[2:0] = 3'b000;
      14'b10000100100111: pixel[2:0] = 3'b000;
      14'b10000100101000: pixel[2:0] = 3'b000;
      14'b10000100101001: pixel[2:0] = 3'b000;
      14'b10000100101010: pixel[2:0] = 3'b000;
      14'b10000100101011: pixel[2:0] = 3'b000;
      14'b10000100101100: pixel[2:0] = 3'b000;
      14'b10000100101101: pixel[2:0] = 3'b000;
      14'b10000100101110: pixel[2:0] = 3'b000;
      14'b10000100101111: pixel[2:0] = 3'b111;
      14'b10000100110000: pixel[2:0] = 3'b111;
      14'b10000100110001: pixel[2:0] = 3'b111;
      14'b10000100110010: pixel[2:0] = 3'b111;
      14'b10000100110011: pixel[2:0] = 3'b111;
      14'b10000100110100: pixel[2:0] = 3'b111;
      14'b10000100110101: pixel[2:0] = 3'b111;
      14'b10000100110110: pixel[2:0] = 3'b111;
      14'b10000100110111: pixel[2:0] = 3'b111;
      14'b10000100111000: pixel[2:0] = 3'b111;
      14'b10000100111001: pixel[2:0] = 3'b111;
      14'b10000100111010: pixel[2:0] = 3'b111;
      14'b10000100111011: pixel[2:0] = 3'b111;
      14'b10000100111100: pixel[2:0] = 3'b111;
      14'b10000100111101: pixel[2:0] = 3'b111;
      14'b10000100111110: pixel[2:0] = 3'b111;
      14'b10000100111111: pixel[2:0] = 3'b111;
      14'b10000101000000: pixel[2:0] = 3'b111;
      14'b10000101000001: pixel[2:0] = 3'b000;
      14'b10000101000010: pixel[2:0] = 3'b000;
      14'b10000101000011: pixel[2:0] = 3'b000;
      14'b10000101000100: pixel[2:0] = 3'b000;
      14'b10000101000101: pixel[2:0] = 3'b000;
      14'b10000101000110: pixel[2:0] = 3'b000;
      14'b10000101000111: pixel[2:0] = 3'b000;
      14'b10000101001000: pixel[2:0] = 3'b000;
      14'b10000101001001: pixel[2:0] = 3'b111;
      14'b10000101001010: pixel[2:0] = 3'b111;
      14'b10000101001011: pixel[2:0] = 3'b111;
      14'b10000101001100: pixel[2:0] = 3'b111;
      14'b10000101001101: pixel[2:0] = 3'b111;
      14'b10000101001110: pixel[2:0] = 3'b000;
      14'b10000101001111: pixel[2:0] = 3'b000;
      14'b10000101010000: pixel[2:0] = 3'b000;
      14'b10000101010001: pixel[2:0] = 3'b000;
      14'b10000101010010: pixel[2:0] = 3'b000;
      14'b10000101010011: pixel[2:0] = 3'b000;
      14'b10000101010100: pixel[2:0] = 3'b000;
      14'b10000101010101: pixel[2:0] = 3'b000;
      14'b10000101010110: pixel[2:0] = 3'b000;
      14'b10000101010111: pixel[2:0] = 3'b000;
      14'b10000101011000: pixel[2:0] = 3'b000;
      14'b10000101011001: pixel[2:0] = 3'b000;
      14'b10000101011010: pixel[2:0] = 3'b111;
      14'b10000101011011: pixel[2:0] = 3'b111;
      14'b10000101011100: pixel[2:0] = 3'b111;
      14'b10000101011101: pixel[2:0] = 3'b111;
      14'b10000101011110: pixel[2:0] = 3'b111;
      14'b10000101011111: pixel[2:0] = 3'b000;
      14'b10000101100000: pixel[2:0] = 3'b000;
      14'b10000101100001: pixel[2:0] = 3'b000;
      14'b10000101100010: pixel[2:0] = 3'b000;
      14'b10000101100011: pixel[2:0] = 3'b000;
      14'b10000101100100: pixel[2:0] = 3'b000;
      14'b10000101100101: pixel[2:0] = 3'b000;
      14'b10000101100110: pixel[2:0] = 3'b000;
      14'b10000101100111: pixel[2:0] = 3'b000;
      14'b10000101101000: pixel[2:0] = 3'b000;
      14'b10000101101001: pixel[2:0] = 3'b000;
      14'b10000101101010: pixel[2:0] = 3'b000;
      14'b10000101101011: pixel[2:0] = 3'b000;
      14'b10000101101100: pixel[2:0] = 3'b000;
      14'b10000101101101: pixel[2:0] = 3'b000;
      14'b10000101101110: pixel[2:0] = 3'b000;
      14'b10000101101111: pixel[2:0] = 3'b000;
      14'b10000101110000: pixel[2:0] = 3'b111;
      14'b10000101110001: pixel[2:0] = 3'b111;
      14'b10000101110010: pixel[2:0] = 3'b111;
      14'b10000101110011: pixel[2:0] = 3'b111;
      14'b10000101110100: pixel[2:0] = 3'b111;
      14'b10000101110101: pixel[2:0] = 3'b000;
      14'b10000101110110: pixel[2:0] = 3'b000;
      14'b10000101110111: pixel[2:0] = 3'b000;
      14'b10000101111000: pixel[2:0] = 3'b000;
      14'b10000101111001: pixel[2:0] = 3'b000;
      14'b10000101111010: pixel[2:0] = 3'b000;
      14'b10000101111011: pixel[2:0] = 3'b000;
      14'b10000101111100: pixel[2:0] = 3'b111;
      14'b10000101111101: pixel[2:0] = 3'b111;
      14'b10000101111110: pixel[2:0] = 3'b111;
      14'b10000101111111: pixel[2:0] = 3'b111;
      14'b10000110000000: pixel[2:0] = 3'b111;
      14'b10000110000001: pixel[2:0] = 3'b000;
      14'b10000110000010: pixel[2:0] = 3'b000;
      14'b10000110000011: pixel[2:0] = 3'b000;
      14'b10000110000100: pixel[2:0] = 3'b000;
      14'b10000110000101: pixel[2:0] = 3'b000;
      14'b10000110000110: pixel[2:0] = 3'b000;
      14'b10000110000111: pixel[2:0] = 3'b000;
      14'b10001000000000: pixel[2:0] = 3'b000;
      14'b10001000000001: pixel[2:0] = 3'b000;
      14'b10001000000010: pixel[2:0] = 3'b111;
      14'b10001000000011: pixel[2:0] = 3'b111;
      14'b10001000000100: pixel[2:0] = 3'b111;
      14'b10001000000101: pixel[2:0] = 3'b111;
      14'b10001000000110: pixel[2:0] = 3'b111;
      14'b10001000000111: pixel[2:0] = 3'b000;
      14'b10001000001000: pixel[2:0] = 3'b000;
      14'b10001000001001: pixel[2:0] = 3'b000;
      14'b10001000001010: pixel[2:0] = 3'b000;
      14'b10001000001011: pixel[2:0] = 3'b000;
      14'b10001000001100: pixel[2:0] = 3'b000;
      14'b10001000001101: pixel[2:0] = 3'b000;
      14'b10001000001110: pixel[2:0] = 3'b000;
      14'b10001000001111: pixel[2:0] = 3'b000;
      14'b10001000010000: pixel[2:0] = 3'b000;
      14'b10001000010001: pixel[2:0] = 3'b000;
      14'b10001000010010: pixel[2:0] = 3'b000;
      14'b10001000010011: pixel[2:0] = 3'b000;
      14'b10001000010100: pixel[2:0] = 3'b000;
      14'b10001000010101: pixel[2:0] = 3'b000;
      14'b10001000010110: pixel[2:0] = 3'b000;
      14'b10001000010111: pixel[2:0] = 3'b000;
      14'b10001000011000: pixel[2:0] = 3'b000;
      14'b10001000011001: pixel[2:0] = 3'b111;
      14'b10001000011010: pixel[2:0] = 3'b111;
      14'b10001000011011: pixel[2:0] = 3'b111;
      14'b10001000011100: pixel[2:0] = 3'b111;
      14'b10001000011101: pixel[2:0] = 3'b111;
      14'b10001000011110: pixel[2:0] = 3'b000;
      14'b10001000011111: pixel[2:0] = 3'b000;
      14'b10001000100000: pixel[2:0] = 3'b000;
      14'b10001000100001: pixel[2:0] = 3'b000;
      14'b10001000100010: pixel[2:0] = 3'b000;
      14'b10001000100011: pixel[2:0] = 3'b000;
      14'b10001000100100: pixel[2:0] = 3'b000;
      14'b10001000100101: pixel[2:0] = 3'b000;
      14'b10001000100110: pixel[2:0] = 3'b000;
      14'b10001000100111: pixel[2:0] = 3'b000;
      14'b10001000101000: pixel[2:0] = 3'b000;
      14'b10001000101001: pixel[2:0] = 3'b000;
      14'b10001000101010: pixel[2:0] = 3'b000;
      14'b10001000101011: pixel[2:0] = 3'b000;
      14'b10001000101100: pixel[2:0] = 3'b000;
      14'b10001000101101: pixel[2:0] = 3'b000;
      14'b10001000101110: pixel[2:0] = 3'b000;
      14'b10001000101111: pixel[2:0] = 3'b111;
      14'b10001000110000: pixel[2:0] = 3'b111;
      14'b10001000110001: pixel[2:0] = 3'b111;
      14'b10001000110010: pixel[2:0] = 3'b111;
      14'b10001000110011: pixel[2:0] = 3'b000;
      14'b10001000110100: pixel[2:0] = 3'b000;
      14'b10001000110101: pixel[2:0] = 3'b000;
      14'b10001000110110: pixel[2:0] = 3'b000;
      14'b10001000110111: pixel[2:0] = 3'b000;
      14'b10001000111000: pixel[2:0] = 3'b000;
      14'b10001000111001: pixel[2:0] = 3'b000;
      14'b10001000111010: pixel[2:0] = 3'b000;
      14'b10001000111011: pixel[2:0] = 3'b000;
      14'b10001000111100: pixel[2:0] = 3'b111;
      14'b10001000111101: pixel[2:0] = 3'b111;
      14'b10001000111110: pixel[2:0] = 3'b111;
      14'b10001000111111: pixel[2:0] = 3'b111;
      14'b10001001000000: pixel[2:0] = 3'b111;
      14'b10001001000001: pixel[2:0] = 3'b000;
      14'b10001001000010: pixel[2:0] = 3'b000;
      14'b10001001000011: pixel[2:0] = 3'b000;
      14'b10001001000100: pixel[2:0] = 3'b000;
      14'b10001001000101: pixel[2:0] = 3'b000;
      14'b10001001000110: pixel[2:0] = 3'b000;
      14'b10001001000111: pixel[2:0] = 3'b000;
      14'b10001001001000: pixel[2:0] = 3'b000;
      14'b10001001001001: pixel[2:0] = 3'b111;
      14'b10001001001010: pixel[2:0] = 3'b111;
      14'b10001001001011: pixel[2:0] = 3'b111;
      14'b10001001001100: pixel[2:0] = 3'b111;
      14'b10001001001101: pixel[2:0] = 3'b111;
      14'b10001001001110: pixel[2:0] = 3'b000;
      14'b10001001001111: pixel[2:0] = 3'b000;
      14'b10001001010000: pixel[2:0] = 3'b000;
      14'b10001001010001: pixel[2:0] = 3'b000;
      14'b10001001010010: pixel[2:0] = 3'b000;
      14'b10001001010011: pixel[2:0] = 3'b000;
      14'b10001001010100: pixel[2:0] = 3'b000;
      14'b10001001010101: pixel[2:0] = 3'b000;
      14'b10001001010110: pixel[2:0] = 3'b000;
      14'b10001001010111: pixel[2:0] = 3'b000;
      14'b10001001011000: pixel[2:0] = 3'b000;
      14'b10001001011001: pixel[2:0] = 3'b000;
      14'b10001001011010: pixel[2:0] = 3'b111;
      14'b10001001011011: pixel[2:0] = 3'b111;
      14'b10001001011100: pixel[2:0] = 3'b111;
      14'b10001001011101: pixel[2:0] = 3'b111;
      14'b10001001011110: pixel[2:0] = 3'b111;
      14'b10001001011111: pixel[2:0] = 3'b000;
      14'b10001001100000: pixel[2:0] = 3'b000;
      14'b10001001100001: pixel[2:0] = 3'b000;
      14'b10001001100010: pixel[2:0] = 3'b000;
      14'b10001001100011: pixel[2:0] = 3'b000;
      14'b10001001100100: pixel[2:0] = 3'b000;
      14'b10001001100101: pixel[2:0] = 3'b000;
      14'b10001001100110: pixel[2:0] = 3'b000;
      14'b10001001100111: pixel[2:0] = 3'b000;
      14'b10001001101000: pixel[2:0] = 3'b000;
      14'b10001001101001: pixel[2:0] = 3'b000;
      14'b10001001101010: pixel[2:0] = 3'b000;
      14'b10001001101011: pixel[2:0] = 3'b000;
      14'b10001001101100: pixel[2:0] = 3'b000;
      14'b10001001101101: pixel[2:0] = 3'b000;
      14'b10001001101110: pixel[2:0] = 3'b000;
      14'b10001001101111: pixel[2:0] = 3'b000;
      14'b10001001110000: pixel[2:0] = 3'b111;
      14'b10001001110001: pixel[2:0] = 3'b111;
      14'b10001001110010: pixel[2:0] = 3'b111;
      14'b10001001110011: pixel[2:0] = 3'b111;
      14'b10001001110100: pixel[2:0] = 3'b111;
      14'b10001001110101: pixel[2:0] = 3'b000;
      14'b10001001110110: pixel[2:0] = 3'b000;
      14'b10001001110111: pixel[2:0] = 3'b000;
      14'b10001001111000: pixel[2:0] = 3'b000;
      14'b10001001111001: pixel[2:0] = 3'b000;
      14'b10001001111010: pixel[2:0] = 3'b000;
      14'b10001001111011: pixel[2:0] = 3'b000;
      14'b10001001111100: pixel[2:0] = 3'b000;
      14'b10001001111101: pixel[2:0] = 3'b111;
      14'b10001001111110: pixel[2:0] = 3'b111;
      14'b10001001111111: pixel[2:0] = 3'b111;
      14'b10001010000000: pixel[2:0] = 3'b111;
      14'b10001010000001: pixel[2:0] = 3'b111;
      14'b10001010000010: pixel[2:0] = 3'b000;
      14'b10001010000011: pixel[2:0] = 3'b000;
      14'b10001010000100: pixel[2:0] = 3'b000;
      14'b10001010000101: pixel[2:0] = 3'b000;
      14'b10001010000110: pixel[2:0] = 3'b000;
      14'b10001010000111: pixel[2:0] = 3'b000;
      14'b10001100000000: pixel[2:0] = 3'b000;
      14'b10001100000001: pixel[2:0] = 3'b000;
      14'b10001100000010: pixel[2:0] = 3'b111;
      14'b10001100000011: pixel[2:0] = 3'b111;
      14'b10001100000100: pixel[2:0] = 3'b111;
      14'b10001100000101: pixel[2:0] = 3'b111;
      14'b10001100000110: pixel[2:0] = 3'b111;
      14'b10001100000111: pixel[2:0] = 3'b000;
      14'b10001100001000: pixel[2:0] = 3'b000;
      14'b10001100001001: pixel[2:0] = 3'b000;
      14'b10001100001010: pixel[2:0] = 3'b000;
      14'b10001100001011: pixel[2:0] = 3'b000;
      14'b10001100001100: pixel[2:0] = 3'b000;
      14'b10001100001101: pixel[2:0] = 3'b000;
      14'b10001100001110: pixel[2:0] = 3'b000;
      14'b10001100001111: pixel[2:0] = 3'b000;
      14'b10001100010000: pixel[2:0] = 3'b000;
      14'b10001100010001: pixel[2:0] = 3'b000;
      14'b10001100010010: pixel[2:0] = 3'b000;
      14'b10001100010011: pixel[2:0] = 3'b000;
      14'b10001100010100: pixel[2:0] = 3'b000;
      14'b10001100010101: pixel[2:0] = 3'b000;
      14'b10001100010110: pixel[2:0] = 3'b000;
      14'b10001100010111: pixel[2:0] = 3'b000;
      14'b10001100011000: pixel[2:0] = 3'b000;
      14'b10001100011001: pixel[2:0] = 3'b111;
      14'b10001100011010: pixel[2:0] = 3'b111;
      14'b10001100011011: pixel[2:0] = 3'b111;
      14'b10001100011100: pixel[2:0] = 3'b111;
      14'b10001100011101: pixel[2:0] = 3'b111;
      14'b10001100011110: pixel[2:0] = 3'b000;
      14'b10001100011111: pixel[2:0] = 3'b000;
      14'b10001100100000: pixel[2:0] = 3'b000;
      14'b10001100100001: pixel[2:0] = 3'b000;
      14'b10001100100010: pixel[2:0] = 3'b000;
      14'b10001100100011: pixel[2:0] = 3'b000;
      14'b10001100100100: pixel[2:0] = 3'b000;
      14'b10001100100101: pixel[2:0] = 3'b000;
      14'b10001100100110: pixel[2:0] = 3'b000;
      14'b10001100100111: pixel[2:0] = 3'b000;
      14'b10001100101000: pixel[2:0] = 3'b000;
      14'b10001100101001: pixel[2:0] = 3'b000;
      14'b10001100101010: pixel[2:0] = 3'b000;
      14'b10001100101011: pixel[2:0] = 3'b000;
      14'b10001100101100: pixel[2:0] = 3'b000;
      14'b10001100101101: pixel[2:0] = 3'b000;
      14'b10001100101110: pixel[2:0] = 3'b111;
      14'b10001100101111: pixel[2:0] = 3'b111;
      14'b10001100110000: pixel[2:0] = 3'b111;
      14'b10001100110001: pixel[2:0] = 3'b111;
      14'b10001100110010: pixel[2:0] = 3'b111;
      14'b10001100110011: pixel[2:0] = 3'b000;
      14'b10001100110100: pixel[2:0] = 3'b000;
      14'b10001100110101: pixel[2:0] = 3'b000;
      14'b10001100110110: pixel[2:0] = 3'b000;
      14'b10001100110111: pixel[2:0] = 3'b000;
      14'b10001100111000: pixel[2:0] = 3'b000;
      14'b10001100111001: pixel[2:0] = 3'b000;
      14'b10001100111010: pixel[2:0] = 3'b000;
      14'b10001100111011: pixel[2:0] = 3'b000;
      14'b10001100111100: pixel[2:0] = 3'b000;
      14'b10001100111101: pixel[2:0] = 3'b111;
      14'b10001100111110: pixel[2:0] = 3'b111;
      14'b10001100111111: pixel[2:0] = 3'b111;
      14'b10001101000000: pixel[2:0] = 3'b111;
      14'b10001101000001: pixel[2:0] = 3'b000;
      14'b10001101000010: pixel[2:0] = 3'b000;
      14'b10001101000011: pixel[2:0] = 3'b000;
      14'b10001101000100: pixel[2:0] = 3'b000;
      14'b10001101000101: pixel[2:0] = 3'b000;
      14'b10001101000110: pixel[2:0] = 3'b000;
      14'b10001101000111: pixel[2:0] = 3'b000;
      14'b10001101001000: pixel[2:0] = 3'b000;
      14'b10001101001001: pixel[2:0] = 3'b111;
      14'b10001101001010: pixel[2:0] = 3'b111;
      14'b10001101001011: pixel[2:0] = 3'b111;
      14'b10001101001100: pixel[2:0] = 3'b111;
      14'b10001101001101: pixel[2:0] = 3'b111;
      14'b10001101001110: pixel[2:0] = 3'b000;
      14'b10001101001111: pixel[2:0] = 3'b000;
      14'b10001101010000: pixel[2:0] = 3'b000;
      14'b10001101010001: pixel[2:0] = 3'b000;
      14'b10001101010010: pixel[2:0] = 3'b000;
      14'b10001101010011: pixel[2:0] = 3'b000;
      14'b10001101010100: pixel[2:0] = 3'b000;
      14'b10001101010101: pixel[2:0] = 3'b000;
      14'b10001101010110: pixel[2:0] = 3'b000;
      14'b10001101010111: pixel[2:0] = 3'b000;
      14'b10001101011000: pixel[2:0] = 3'b000;
      14'b10001101011001: pixel[2:0] = 3'b000;
      14'b10001101011010: pixel[2:0] = 3'b111;
      14'b10001101011011: pixel[2:0] = 3'b111;
      14'b10001101011100: pixel[2:0] = 3'b111;
      14'b10001101011101: pixel[2:0] = 3'b111;
      14'b10001101011110: pixel[2:0] = 3'b111;
      14'b10001101011111: pixel[2:0] = 3'b000;
      14'b10001101100000: pixel[2:0] = 3'b000;
      14'b10001101100001: pixel[2:0] = 3'b000;
      14'b10001101100010: pixel[2:0] = 3'b000;
      14'b10001101100011: pixel[2:0] = 3'b000;
      14'b10001101100100: pixel[2:0] = 3'b000;
      14'b10001101100101: pixel[2:0] = 3'b000;
      14'b10001101100110: pixel[2:0] = 3'b000;
      14'b10001101100111: pixel[2:0] = 3'b000;
      14'b10001101101000: pixel[2:0] = 3'b000;
      14'b10001101101001: pixel[2:0] = 3'b000;
      14'b10001101101010: pixel[2:0] = 3'b000;
      14'b10001101101011: pixel[2:0] = 3'b000;
      14'b10001101101100: pixel[2:0] = 3'b000;
      14'b10001101101101: pixel[2:0] = 3'b000;
      14'b10001101101110: pixel[2:0] = 3'b000;
      14'b10001101101111: pixel[2:0] = 3'b000;
      14'b10001101110000: pixel[2:0] = 3'b111;
      14'b10001101110001: pixel[2:0] = 3'b111;
      14'b10001101110010: pixel[2:0] = 3'b111;
      14'b10001101110011: pixel[2:0] = 3'b111;
      14'b10001101110100: pixel[2:0] = 3'b111;
      14'b10001101110101: pixel[2:0] = 3'b000;
      14'b10001101110110: pixel[2:0] = 3'b000;
      14'b10001101110111: pixel[2:0] = 3'b000;
      14'b10001101111000: pixel[2:0] = 3'b000;
      14'b10001101111001: pixel[2:0] = 3'b000;
      14'b10001101111010: pixel[2:0] = 3'b000;
      14'b10001101111011: pixel[2:0] = 3'b000;
      14'b10001101111100: pixel[2:0] = 3'b000;
      14'b10001101111101: pixel[2:0] = 3'b111;
      14'b10001101111110: pixel[2:0] = 3'b111;
      14'b10001101111111: pixel[2:0] = 3'b111;
      14'b10001110000000: pixel[2:0] = 3'b111;
      14'b10001110000001: pixel[2:0] = 3'b111;
      14'b10001110000010: pixel[2:0] = 3'b000;
      14'b10001110000011: pixel[2:0] = 3'b000;
      14'b10001110000100: pixel[2:0] = 3'b000;
      14'b10001110000101: pixel[2:0] = 3'b000;
      14'b10001110000110: pixel[2:0] = 3'b000;
      14'b10001110000111: pixel[2:0] = 3'b000;
      14'b10010000000000: pixel[2:0] = 3'b000;
      14'b10010000000001: pixel[2:0] = 3'b000;
      14'b10010000000010: pixel[2:0] = 3'b111;
      14'b10010000000011: pixel[2:0] = 3'b111;
      14'b10010000000100: pixel[2:0] = 3'b111;
      14'b10010000000101: pixel[2:0] = 3'b111;
      14'b10010000000110: pixel[2:0] = 3'b111;
      14'b10010000000111: pixel[2:0] = 3'b000;
      14'b10010000001000: pixel[2:0] = 3'b000;
      14'b10010000001001: pixel[2:0] = 3'b000;
      14'b10010000001010: pixel[2:0] = 3'b000;
      14'b10010000001011: pixel[2:0] = 3'b000;
      14'b10010000001100: pixel[2:0] = 3'b000;
      14'b10010000001101: pixel[2:0] = 3'b000;
      14'b10010000001110: pixel[2:0] = 3'b000;
      14'b10010000001111: pixel[2:0] = 3'b000;
      14'b10010000010000: pixel[2:0] = 3'b000;
      14'b10010000010001: pixel[2:0] = 3'b000;
      14'b10010000010010: pixel[2:0] = 3'b000;
      14'b10010000010011: pixel[2:0] = 3'b000;
      14'b10010000010100: pixel[2:0] = 3'b000;
      14'b10010000010101: pixel[2:0] = 3'b000;
      14'b10010000010110: pixel[2:0] = 3'b000;
      14'b10010000010111: pixel[2:0] = 3'b000;
      14'b10010000011000: pixel[2:0] = 3'b000;
      14'b10010000011001: pixel[2:0] = 3'b111;
      14'b10010000011010: pixel[2:0] = 3'b111;
      14'b10010000011011: pixel[2:0] = 3'b111;
      14'b10010000011100: pixel[2:0] = 3'b111;
      14'b10010000011101: pixel[2:0] = 3'b111;
      14'b10010000011110: pixel[2:0] = 3'b000;
      14'b10010000011111: pixel[2:0] = 3'b000;
      14'b10010000100000: pixel[2:0] = 3'b000;
      14'b10010000100001: pixel[2:0] = 3'b000;
      14'b10010000100010: pixel[2:0] = 3'b000;
      14'b10010000100011: pixel[2:0] = 3'b000;
      14'b10010000100100: pixel[2:0] = 3'b000;
      14'b10010000100101: pixel[2:0] = 3'b000;
      14'b10010000100110: pixel[2:0] = 3'b000;
      14'b10010000100111: pixel[2:0] = 3'b000;
      14'b10010000101000: pixel[2:0] = 3'b000;
      14'b10010000101001: pixel[2:0] = 3'b000;
      14'b10010000101010: pixel[2:0] = 3'b000;
      14'b10010000101011: pixel[2:0] = 3'b000;
      14'b10010000101100: pixel[2:0] = 3'b000;
      14'b10010000101101: pixel[2:0] = 3'b000;
      14'b10010000101110: pixel[2:0] = 3'b111;
      14'b10010000101111: pixel[2:0] = 3'b111;
      14'b10010000110000: pixel[2:0] = 3'b111;
      14'b10010000110001: pixel[2:0] = 3'b111;
      14'b10010000110010: pixel[2:0] = 3'b111;
      14'b10010000110011: pixel[2:0] = 3'b000;
      14'b10010000110100: pixel[2:0] = 3'b000;
      14'b10010000110101: pixel[2:0] = 3'b000;
      14'b10010000110110: pixel[2:0] = 3'b000;
      14'b10010000110111: pixel[2:0] = 3'b000;
      14'b10010000111000: pixel[2:0] = 3'b000;
      14'b10010000111001: pixel[2:0] = 3'b000;
      14'b10010000111010: pixel[2:0] = 3'b000;
      14'b10010000111011: pixel[2:0] = 3'b000;
      14'b10010000111100: pixel[2:0] = 3'b000;
      14'b10010000111101: pixel[2:0] = 3'b111;
      14'b10010000111110: pixel[2:0] = 3'b111;
      14'b10010000111111: pixel[2:0] = 3'b111;
      14'b10010001000000: pixel[2:0] = 3'b111;
      14'b10010001000001: pixel[2:0] = 3'b111;
      14'b10010001000010: pixel[2:0] = 3'b000;
      14'b10010001000011: pixel[2:0] = 3'b000;
      14'b10010001000100: pixel[2:0] = 3'b000;
      14'b10010001000101: pixel[2:0] = 3'b000;
      14'b10010001000110: pixel[2:0] = 3'b000;
      14'b10010001000111: pixel[2:0] = 3'b000;
      14'b10010001001000: pixel[2:0] = 3'b000;
      14'b10010001001001: pixel[2:0] = 3'b111;
      14'b10010001001010: pixel[2:0] = 3'b111;
      14'b10010001001011: pixel[2:0] = 3'b111;
      14'b10010001001100: pixel[2:0] = 3'b111;
      14'b10010001001101: pixel[2:0] = 3'b111;
      14'b10010001001110: pixel[2:0] = 3'b000;
      14'b10010001001111: pixel[2:0] = 3'b000;
      14'b10010001010000: pixel[2:0] = 3'b000;
      14'b10010001010001: pixel[2:0] = 3'b000;
      14'b10010001010010: pixel[2:0] = 3'b000;
      14'b10010001010011: pixel[2:0] = 3'b000;
      14'b10010001010100: pixel[2:0] = 3'b000;
      14'b10010001010101: pixel[2:0] = 3'b000;
      14'b10010001010110: pixel[2:0] = 3'b000;
      14'b10010001010111: pixel[2:0] = 3'b000;
      14'b10010001011000: pixel[2:0] = 3'b000;
      14'b10010001011001: pixel[2:0] = 3'b000;
      14'b10010001011010: pixel[2:0] = 3'b111;
      14'b10010001011011: pixel[2:0] = 3'b111;
      14'b10010001011100: pixel[2:0] = 3'b111;
      14'b10010001011101: pixel[2:0] = 3'b111;
      14'b10010001011110: pixel[2:0] = 3'b111;
      14'b10010001011111: pixel[2:0] = 3'b000;
      14'b10010001100000: pixel[2:0] = 3'b000;
      14'b10010001100001: pixel[2:0] = 3'b000;
      14'b10010001100010: pixel[2:0] = 3'b000;
      14'b10010001100011: pixel[2:0] = 3'b000;
      14'b10010001100100: pixel[2:0] = 3'b000;
      14'b10010001100101: pixel[2:0] = 3'b000;
      14'b10010001100110: pixel[2:0] = 3'b000;
      14'b10010001100111: pixel[2:0] = 3'b000;
      14'b10010001101000: pixel[2:0] = 3'b000;
      14'b10010001101001: pixel[2:0] = 3'b000;
      14'b10010001101010: pixel[2:0] = 3'b000;
      14'b10010001101011: pixel[2:0] = 3'b000;
      14'b10010001101100: pixel[2:0] = 3'b000;
      14'b10010001101101: pixel[2:0] = 3'b000;
      14'b10010001101110: pixel[2:0] = 3'b000;
      14'b10010001101111: pixel[2:0] = 3'b000;
      14'b10010001110000: pixel[2:0] = 3'b111;
      14'b10010001110001: pixel[2:0] = 3'b111;
      14'b10010001110010: pixel[2:0] = 3'b111;
      14'b10010001110011: pixel[2:0] = 3'b111;
      14'b10010001110100: pixel[2:0] = 3'b111;
      14'b10010001110101: pixel[2:0] = 3'b000;
      14'b10010001110110: pixel[2:0] = 3'b000;
      14'b10010001110111: pixel[2:0] = 3'b000;
      14'b10010001111000: pixel[2:0] = 3'b000;
      14'b10010001111001: pixel[2:0] = 3'b000;
      14'b10010001111010: pixel[2:0] = 3'b000;
      14'b10010001111011: pixel[2:0] = 3'b000;
      14'b10010001111100: pixel[2:0] = 3'b000;
      14'b10010001111101: pixel[2:0] = 3'b111;
      14'b10010001111110: pixel[2:0] = 3'b111;
      14'b10010001111111: pixel[2:0] = 3'b111;
      14'b10010010000000: pixel[2:0] = 3'b111;
      14'b10010010000001: pixel[2:0] = 3'b111;
      14'b10010010000010: pixel[2:0] = 3'b000;
      14'b10010010000011: pixel[2:0] = 3'b000;
      14'b10010010000100: pixel[2:0] = 3'b000;
      14'b10010010000101: pixel[2:0] = 3'b000;
      14'b10010010000110: pixel[2:0] = 3'b000;
      14'b10010010000111: pixel[2:0] = 3'b000;
      14'b10010100000000: pixel[2:0] = 3'b000;
      14'b10010100000001: pixel[2:0] = 3'b000;
      14'b10010100000010: pixel[2:0] = 3'b111;
      14'b10010100000011: pixel[2:0] = 3'b111;
      14'b10010100000100: pixel[2:0] = 3'b111;
      14'b10010100000101: pixel[2:0] = 3'b111;
      14'b10010100000110: pixel[2:0] = 3'b111;
      14'b10010100000111: pixel[2:0] = 3'b000;
      14'b10010100001000: pixel[2:0] = 3'b000;
      14'b10010100001001: pixel[2:0] = 3'b000;
      14'b10010100001010: pixel[2:0] = 3'b000;
      14'b10010100001011: pixel[2:0] = 3'b000;
      14'b10010100001100: pixel[2:0] = 3'b000;
      14'b10010100001101: pixel[2:0] = 3'b000;
      14'b10010100001110: pixel[2:0] = 3'b000;
      14'b10010100001111: pixel[2:0] = 3'b000;
      14'b10010100010000: pixel[2:0] = 3'b000;
      14'b10010100010001: pixel[2:0] = 3'b000;
      14'b10010100010010: pixel[2:0] = 3'b000;
      14'b10010100010011: pixel[2:0] = 3'b000;
      14'b10010100010100: pixel[2:0] = 3'b000;
      14'b10010100010101: pixel[2:0] = 3'b000;
      14'b10010100010110: pixel[2:0] = 3'b000;
      14'b10010100010111: pixel[2:0] = 3'b000;
      14'b10010100011000: pixel[2:0] = 3'b000;
      14'b10010100011001: pixel[2:0] = 3'b111;
      14'b10010100011010: pixel[2:0] = 3'b111;
      14'b10010100011011: pixel[2:0] = 3'b111;
      14'b10010100011100: pixel[2:0] = 3'b111;
      14'b10010100011101: pixel[2:0] = 3'b111;
      14'b10010100011110: pixel[2:0] = 3'b111;
      14'b10010100011111: pixel[2:0] = 3'b111;
      14'b10010100100000: pixel[2:0] = 3'b111;
      14'b10010100100001: pixel[2:0] = 3'b111;
      14'b10010100100010: pixel[2:0] = 3'b111;
      14'b10010100100011: pixel[2:0] = 3'b111;
      14'b10010100100100: pixel[2:0] = 3'b111;
      14'b10010100100101: pixel[2:0] = 3'b111;
      14'b10010100100110: pixel[2:0] = 3'b111;
      14'b10010100100111: pixel[2:0] = 3'b111;
      14'b10010100101000: pixel[2:0] = 3'b111;
      14'b10010100101001: pixel[2:0] = 3'b111;
      14'b10010100101010: pixel[2:0] = 3'b000;
      14'b10010100101011: pixel[2:0] = 3'b000;
      14'b10010100101100: pixel[2:0] = 3'b000;
      14'b10010100101101: pixel[2:0] = 3'b000;
      14'b10010100101110: pixel[2:0] = 3'b111;
      14'b10010100101111: pixel[2:0] = 3'b111;
      14'b10010100110000: pixel[2:0] = 3'b111;
      14'b10010100110001: pixel[2:0] = 3'b111;
      14'b10010100110010: pixel[2:0] = 3'b111;
      14'b10010100110011: pixel[2:0] = 3'b000;
      14'b10010100110100: pixel[2:0] = 3'b000;
      14'b10010100110101: pixel[2:0] = 3'b000;
      14'b10010100110110: pixel[2:0] = 3'b000;
      14'b10010100110111: pixel[2:0] = 3'b000;
      14'b10010100111000: pixel[2:0] = 3'b000;
      14'b10010100111001: pixel[2:0] = 3'b000;
      14'b10010100111010: pixel[2:0] = 3'b000;
      14'b10010100111011: pixel[2:0] = 3'b000;
      14'b10010100111100: pixel[2:0] = 3'b000;
      14'b10010100111101: pixel[2:0] = 3'b111;
      14'b10010100111110: pixel[2:0] = 3'b111;
      14'b10010100111111: pixel[2:0] = 3'b111;
      14'b10010101000000: pixel[2:0] = 3'b111;
      14'b10010101000001: pixel[2:0] = 3'b111;
      14'b10010101000010: pixel[2:0] = 3'b000;
      14'b10010101000011: pixel[2:0] = 3'b000;
      14'b10010101000100: pixel[2:0] = 3'b000;
      14'b10010101000101: pixel[2:0] = 3'b000;
      14'b10010101000110: pixel[2:0] = 3'b000;
      14'b10010101000111: pixel[2:0] = 3'b000;
      14'b10010101001000: pixel[2:0] = 3'b000;
      14'b10010101001001: pixel[2:0] = 3'b111;
      14'b10010101001010: pixel[2:0] = 3'b111;
      14'b10010101001011: pixel[2:0] = 3'b111;
      14'b10010101001100: pixel[2:0] = 3'b111;
      14'b10010101001101: pixel[2:0] = 3'b111;
      14'b10010101001110: pixel[2:0] = 3'b000;
      14'b10010101001111: pixel[2:0] = 3'b000;
      14'b10010101010000: pixel[2:0] = 3'b000;
      14'b10010101010001: pixel[2:0] = 3'b000;
      14'b10010101010010: pixel[2:0] = 3'b000;
      14'b10010101010011: pixel[2:0] = 3'b000;
      14'b10010101010100: pixel[2:0] = 3'b000;
      14'b10010101010101: pixel[2:0] = 3'b000;
      14'b10010101010110: pixel[2:0] = 3'b000;
      14'b10010101010111: pixel[2:0] = 3'b000;
      14'b10010101011000: pixel[2:0] = 3'b000;
      14'b10010101011001: pixel[2:0] = 3'b000;
      14'b10010101011010: pixel[2:0] = 3'b111;
      14'b10010101011011: pixel[2:0] = 3'b111;
      14'b10010101011100: pixel[2:0] = 3'b111;
      14'b10010101011101: pixel[2:0] = 3'b111;
      14'b10010101011110: pixel[2:0] = 3'b111;
      14'b10010101011111: pixel[2:0] = 3'b111;
      14'b10010101100000: pixel[2:0] = 3'b111;
      14'b10010101100001: pixel[2:0] = 3'b111;
      14'b10010101100010: pixel[2:0] = 3'b111;
      14'b10010101100011: pixel[2:0] = 3'b111;
      14'b10010101100100: pixel[2:0] = 3'b111;
      14'b10010101100101: pixel[2:0] = 3'b111;
      14'b10010101100110: pixel[2:0] = 3'b111;
      14'b10010101100111: pixel[2:0] = 3'b111;
      14'b10010101101000: pixel[2:0] = 3'b111;
      14'b10010101101001: pixel[2:0] = 3'b111;
      14'b10010101101010: pixel[2:0] = 3'b111;
      14'b10010101101011: pixel[2:0] = 3'b000;
      14'b10010101101100: pixel[2:0] = 3'b000;
      14'b10010101101101: pixel[2:0] = 3'b000;
      14'b10010101101110: pixel[2:0] = 3'b000;
      14'b10010101101111: pixel[2:0] = 3'b000;
      14'b10010101110000: pixel[2:0] = 3'b111;
      14'b10010101110001: pixel[2:0] = 3'b111;
      14'b10010101110010: pixel[2:0] = 3'b111;
      14'b10010101110011: pixel[2:0] = 3'b111;
      14'b10010101110100: pixel[2:0] = 3'b111;
      14'b10010101110101: pixel[2:0] = 3'b000;
      14'b10010101110110: pixel[2:0] = 3'b000;
      14'b10010101110111: pixel[2:0] = 3'b000;
      14'b10010101111000: pixel[2:0] = 3'b000;
      14'b10010101111001: pixel[2:0] = 3'b000;
      14'b10010101111010: pixel[2:0] = 3'b000;
      14'b10010101111011: pixel[2:0] = 3'b000;
      14'b10010101111100: pixel[2:0] = 3'b000;
      14'b10010101111101: pixel[2:0] = 3'b111;
      14'b10010101111110: pixel[2:0] = 3'b111;
      14'b10010101111111: pixel[2:0] = 3'b111;
      14'b10010110000000: pixel[2:0] = 3'b111;
      14'b10010110000001: pixel[2:0] = 3'b111;
      14'b10010110000010: pixel[2:0] = 3'b111;
      14'b10010110000011: pixel[2:0] = 3'b000;
      14'b10010110000100: pixel[2:0] = 3'b000;
      14'b10010110000101: pixel[2:0] = 3'b000;
      14'b10010110000110: pixel[2:0] = 3'b000;
      14'b10010110000111: pixel[2:0] = 3'b000;
      14'b10011000000000: pixel[2:0] = 3'b000;
      14'b10011000000001: pixel[2:0] = 3'b000;
      14'b10011000000010: pixel[2:0] = 3'b111;
      14'b10011000000011: pixel[2:0] = 3'b111;
      14'b10011000000100: pixel[2:0] = 3'b111;
      14'b10011000000101: pixel[2:0] = 3'b111;
      14'b10011000000110: pixel[2:0] = 3'b111;
      14'b10011000000111: pixel[2:0] = 3'b000;
      14'b10011000001000: pixel[2:0] = 3'b000;
      14'b10011000001001: pixel[2:0] = 3'b000;
      14'b10011000001010: pixel[2:0] = 3'b000;
      14'b10011000001011: pixel[2:0] = 3'b000;
      14'b10011000001100: pixel[2:0] = 3'b000;
      14'b10011000001101: pixel[2:0] = 3'b000;
      14'b10011000001110: pixel[2:0] = 3'b000;
      14'b10011000001111: pixel[2:0] = 3'b000;
      14'b10011000010000: pixel[2:0] = 3'b000;
      14'b10011000010001: pixel[2:0] = 3'b000;
      14'b10011000010010: pixel[2:0] = 3'b000;
      14'b10011000010011: pixel[2:0] = 3'b000;
      14'b10011000010100: pixel[2:0] = 3'b000;
      14'b10011000010101: pixel[2:0] = 3'b000;
      14'b10011000010110: pixel[2:0] = 3'b000;
      14'b10011000010111: pixel[2:0] = 3'b000;
      14'b10011000011000: pixel[2:0] = 3'b000;
      14'b10011000011001: pixel[2:0] = 3'b111;
      14'b10011000011010: pixel[2:0] = 3'b111;
      14'b10011000011011: pixel[2:0] = 3'b111;
      14'b10011000011100: pixel[2:0] = 3'b111;
      14'b10011000011101: pixel[2:0] = 3'b111;
      14'b10011000011110: pixel[2:0] = 3'b111;
      14'b10011000011111: pixel[2:0] = 3'b111;
      14'b10011000100000: pixel[2:0] = 3'b111;
      14'b10011000100001: pixel[2:0] = 3'b111;
      14'b10011000100010: pixel[2:0] = 3'b111;
      14'b10011000100011: pixel[2:0] = 3'b111;
      14'b10011000100100: pixel[2:0] = 3'b111;
      14'b10011000100101: pixel[2:0] = 3'b111;
      14'b10011000100110: pixel[2:0] = 3'b111;
      14'b10011000100111: pixel[2:0] = 3'b111;
      14'b10011000101000: pixel[2:0] = 3'b111;
      14'b10011000101001: pixel[2:0] = 3'b111;
      14'b10011000101010: pixel[2:0] = 3'b000;
      14'b10011000101011: pixel[2:0] = 3'b000;
      14'b10011000101100: pixel[2:0] = 3'b000;
      14'b10011000101101: pixel[2:0] = 3'b000;
      14'b10011000101110: pixel[2:0] = 3'b111;
      14'b10011000101111: pixel[2:0] = 3'b111;
      14'b10011000110000: pixel[2:0] = 3'b111;
      14'b10011000110001: pixel[2:0] = 3'b111;
      14'b10011000110010: pixel[2:0] = 3'b000;
      14'b10011000110011: pixel[2:0] = 3'b000;
      14'b10011000110100: pixel[2:0] = 3'b000;
      14'b10011000110101: pixel[2:0] = 3'b000;
      14'b10011000110110: pixel[2:0] = 3'b000;
      14'b10011000110111: pixel[2:0] = 3'b000;
      14'b10011000111000: pixel[2:0] = 3'b000;
      14'b10011000111001: pixel[2:0] = 3'b000;
      14'b10011000111010: pixel[2:0] = 3'b000;
      14'b10011000111011: pixel[2:0] = 3'b000;
      14'b10011000111100: pixel[2:0] = 3'b000;
      14'b10011000111101: pixel[2:0] = 3'b111;
      14'b10011000111110: pixel[2:0] = 3'b111;
      14'b10011000111111: pixel[2:0] = 3'b111;
      14'b10011001000000: pixel[2:0] = 3'b111;
      14'b10011001000001: pixel[2:0] = 3'b111;
      14'b10011001000010: pixel[2:0] = 3'b000;
      14'b10011001000011: pixel[2:0] = 3'b000;
      14'b10011001000100: pixel[2:0] = 3'b000;
      14'b10011001000101: pixel[2:0] = 3'b000;
      14'b10011001000110: pixel[2:0] = 3'b000;
      14'b10011001000111: pixel[2:0] = 3'b000;
      14'b10011001001000: pixel[2:0] = 3'b000;
      14'b10011001001001: pixel[2:0] = 3'b111;
      14'b10011001001010: pixel[2:0] = 3'b111;
      14'b10011001001011: pixel[2:0] = 3'b111;
      14'b10011001001100: pixel[2:0] = 3'b111;
      14'b10011001001101: pixel[2:0] = 3'b111;
      14'b10011001001110: pixel[2:0] = 3'b000;
      14'b10011001001111: pixel[2:0] = 3'b000;
      14'b10011001010000: pixel[2:0] = 3'b000;
      14'b10011001010001: pixel[2:0] = 3'b000;
      14'b10011001010010: pixel[2:0] = 3'b000;
      14'b10011001010011: pixel[2:0] = 3'b000;
      14'b10011001010100: pixel[2:0] = 3'b000;
      14'b10011001010101: pixel[2:0] = 3'b000;
      14'b10011001010110: pixel[2:0] = 3'b000;
      14'b10011001010111: pixel[2:0] = 3'b000;
      14'b10011001011000: pixel[2:0] = 3'b000;
      14'b10011001011001: pixel[2:0] = 3'b000;
      14'b10011001011010: pixel[2:0] = 3'b111;
      14'b10011001011011: pixel[2:0] = 3'b111;
      14'b10011001011100: pixel[2:0] = 3'b111;
      14'b10011001011101: pixel[2:0] = 3'b111;
      14'b10011001011110: pixel[2:0] = 3'b111;
      14'b10011001011111: pixel[2:0] = 3'b111;
      14'b10011001100000: pixel[2:0] = 3'b111;
      14'b10011001100001: pixel[2:0] = 3'b111;
      14'b10011001100010: pixel[2:0] = 3'b111;
      14'b10011001100011: pixel[2:0] = 3'b111;
      14'b10011001100100: pixel[2:0] = 3'b111;
      14'b10011001100101: pixel[2:0] = 3'b111;
      14'b10011001100110: pixel[2:0] = 3'b111;
      14'b10011001100111: pixel[2:0] = 3'b111;
      14'b10011001101000: pixel[2:0] = 3'b111;
      14'b10011001101001: pixel[2:0] = 3'b111;
      14'b10011001101010: pixel[2:0] = 3'b111;
      14'b10011001101011: pixel[2:0] = 3'b000;
      14'b10011001101100: pixel[2:0] = 3'b000;
      14'b10011001101101: pixel[2:0] = 3'b000;
      14'b10011001101110: pixel[2:0] = 3'b000;
      14'b10011001101111: pixel[2:0] = 3'b000;
      14'b10011001110000: pixel[2:0] = 3'b111;
      14'b10011001110001: pixel[2:0] = 3'b111;
      14'b10011001110010: pixel[2:0] = 3'b111;
      14'b10011001110011: pixel[2:0] = 3'b111;
      14'b10011001110100: pixel[2:0] = 3'b111;
      14'b10011001110101: pixel[2:0] = 3'b000;
      14'b10011001110110: pixel[2:0] = 3'b000;
      14'b10011001110111: pixel[2:0] = 3'b000;
      14'b10011001111000: pixel[2:0] = 3'b000;
      14'b10011001111001: pixel[2:0] = 3'b000;
      14'b10011001111010: pixel[2:0] = 3'b000;
      14'b10011001111011: pixel[2:0] = 3'b000;
      14'b10011001111100: pixel[2:0] = 3'b000;
      14'b10011001111101: pixel[2:0] = 3'b000;
      14'b10011001111110: pixel[2:0] = 3'b111;
      14'b10011001111111: pixel[2:0] = 3'b111;
      14'b10011010000000: pixel[2:0] = 3'b111;
      14'b10011010000001: pixel[2:0] = 3'b111;
      14'b10011010000010: pixel[2:0] = 3'b111;
      14'b10011010000011: pixel[2:0] = 3'b000;
      14'b10011010000100: pixel[2:0] = 3'b000;
      14'b10011010000101: pixel[2:0] = 3'b000;
      14'b10011010000110: pixel[2:0] = 3'b000;
      14'b10011010000111: pixel[2:0] = 3'b000;
      14'b10011100000000: pixel[2:0] = 3'b000;
      14'b10011100000001: pixel[2:0] = 3'b000;
      14'b10011100000010: pixel[2:0] = 3'b111;
      14'b10011100000011: pixel[2:0] = 3'b111;
      14'b10011100000100: pixel[2:0] = 3'b111;
      14'b10011100000101: pixel[2:0] = 3'b111;
      14'b10011100000110: pixel[2:0] = 3'b111;
      14'b10011100000111: pixel[2:0] = 3'b000;
      14'b10011100001000: pixel[2:0] = 3'b000;
      14'b10011100001001: pixel[2:0] = 3'b000;
      14'b10011100001010: pixel[2:0] = 3'b000;
      14'b10011100001011: pixel[2:0] = 3'b000;
      14'b10011100001100: pixel[2:0] = 3'b000;
      14'b10011100001101: pixel[2:0] = 3'b000;
      14'b10011100001110: pixel[2:0] = 3'b000;
      14'b10011100001111: pixel[2:0] = 3'b000;
      14'b10011100010000: pixel[2:0] = 3'b000;
      14'b10011100010001: pixel[2:0] = 3'b000;
      14'b10011100010010: pixel[2:0] = 3'b000;
      14'b10011100010011: pixel[2:0] = 3'b000;
      14'b10011100010100: pixel[2:0] = 3'b000;
      14'b10011100010101: pixel[2:0] = 3'b000;
      14'b10011100010110: pixel[2:0] = 3'b000;
      14'b10011100010111: pixel[2:0] = 3'b000;
      14'b10011100011000: pixel[2:0] = 3'b000;
      14'b10011100011001: pixel[2:0] = 3'b111;
      14'b10011100011010: pixel[2:0] = 3'b111;
      14'b10011100011011: pixel[2:0] = 3'b111;
      14'b10011100011100: pixel[2:0] = 3'b111;
      14'b10011100011101: pixel[2:0] = 3'b111;
      14'b10011100011110: pixel[2:0] = 3'b111;
      14'b10011100011111: pixel[2:0] = 3'b111;
      14'b10011100100000: pixel[2:0] = 3'b111;
      14'b10011100100001: pixel[2:0] = 3'b111;
      14'b10011100100010: pixel[2:0] = 3'b111;
      14'b10011100100011: pixel[2:0] = 3'b111;
      14'b10011100100100: pixel[2:0] = 3'b111;
      14'b10011100100101: pixel[2:0] = 3'b111;
      14'b10011100100110: pixel[2:0] = 3'b111;
      14'b10011100100111: pixel[2:0] = 3'b111;
      14'b10011100101000: pixel[2:0] = 3'b111;
      14'b10011100101001: pixel[2:0] = 3'b111;
      14'b10011100101010: pixel[2:0] = 3'b000;
      14'b10011100101011: pixel[2:0] = 3'b000;
      14'b10011100101100: pixel[2:0] = 3'b000;
      14'b10011100101101: pixel[2:0] = 3'b111;
      14'b10011100101110: pixel[2:0] = 3'b111;
      14'b10011100101111: pixel[2:0] = 3'b111;
      14'b10011100110000: pixel[2:0] = 3'b111;
      14'b10011100110001: pixel[2:0] = 3'b111;
      14'b10011100110010: pixel[2:0] = 3'b000;
      14'b10011100110011: pixel[2:0] = 3'b000;
      14'b10011100110100: pixel[2:0] = 3'b000;
      14'b10011100110101: pixel[2:0] = 3'b000;
      14'b10011100110110: pixel[2:0] = 3'b000;
      14'b10011100110111: pixel[2:0] = 3'b000;
      14'b10011100111000: pixel[2:0] = 3'b000;
      14'b10011100111001: pixel[2:0] = 3'b000;
      14'b10011100111010: pixel[2:0] = 3'b000;
      14'b10011100111011: pixel[2:0] = 3'b000;
      14'b10011100111100: pixel[2:0] = 3'b000;
      14'b10011100111101: pixel[2:0] = 3'b111;
      14'b10011100111110: pixel[2:0] = 3'b111;
      14'b10011100111111: pixel[2:0] = 3'b111;
      14'b10011101000000: pixel[2:0] = 3'b111;
      14'b10011101000001: pixel[2:0] = 3'b111;
      14'b10011101000010: pixel[2:0] = 3'b000;
      14'b10011101000011: pixel[2:0] = 3'b000;
      14'b10011101000100: pixel[2:0] = 3'b000;
      14'b10011101000101: pixel[2:0] = 3'b000;
      14'b10011101000110: pixel[2:0] = 3'b000;
      14'b10011101000111: pixel[2:0] = 3'b000;
      14'b10011101001000: pixel[2:0] = 3'b000;
      14'b10011101001001: pixel[2:0] = 3'b111;
      14'b10011101001010: pixel[2:0] = 3'b111;
      14'b10011101001011: pixel[2:0] = 3'b111;
      14'b10011101001100: pixel[2:0] = 3'b111;
      14'b10011101001101: pixel[2:0] = 3'b111;
      14'b10011101001110: pixel[2:0] = 3'b000;
      14'b10011101001111: pixel[2:0] = 3'b000;
      14'b10011101010000: pixel[2:0] = 3'b000;
      14'b10011101010001: pixel[2:0] = 3'b000;
      14'b10011101010010: pixel[2:0] = 3'b000;
      14'b10011101010011: pixel[2:0] = 3'b000;
      14'b10011101010100: pixel[2:0] = 3'b000;
      14'b10011101010101: pixel[2:0] = 3'b000;
      14'b10011101010110: pixel[2:0] = 3'b000;
      14'b10011101010111: pixel[2:0] = 3'b000;
      14'b10011101011000: pixel[2:0] = 3'b000;
      14'b10011101011001: pixel[2:0] = 3'b000;
      14'b10011101011010: pixel[2:0] = 3'b111;
      14'b10011101011011: pixel[2:0] = 3'b111;
      14'b10011101011100: pixel[2:0] = 3'b111;
      14'b10011101011101: pixel[2:0] = 3'b111;
      14'b10011101011110: pixel[2:0] = 3'b111;
      14'b10011101011111: pixel[2:0] = 3'b111;
      14'b10011101100000: pixel[2:0] = 3'b111;
      14'b10011101100001: pixel[2:0] = 3'b111;
      14'b10011101100010: pixel[2:0] = 3'b111;
      14'b10011101100011: pixel[2:0] = 3'b111;
      14'b10011101100100: pixel[2:0] = 3'b111;
      14'b10011101100101: pixel[2:0] = 3'b111;
      14'b10011101100110: pixel[2:0] = 3'b111;
      14'b10011101100111: pixel[2:0] = 3'b111;
      14'b10011101101000: pixel[2:0] = 3'b111;
      14'b10011101101001: pixel[2:0] = 3'b111;
      14'b10011101101010: pixel[2:0] = 3'b111;
      14'b10011101101011: pixel[2:0] = 3'b000;
      14'b10011101101100: pixel[2:0] = 3'b000;
      14'b10011101101101: pixel[2:0] = 3'b000;
      14'b10011101101110: pixel[2:0] = 3'b000;
      14'b10011101101111: pixel[2:0] = 3'b000;
      14'b10011101110000: pixel[2:0] = 3'b111;
      14'b10011101110001: pixel[2:0] = 3'b111;
      14'b10011101110010: pixel[2:0] = 3'b111;
      14'b10011101110011: pixel[2:0] = 3'b111;
      14'b10011101110100: pixel[2:0] = 3'b111;
      14'b10011101110101: pixel[2:0] = 3'b000;
      14'b10011101110110: pixel[2:0] = 3'b000;
      14'b10011101110111: pixel[2:0] = 3'b000;
      14'b10011101111000: pixel[2:0] = 3'b000;
      14'b10011101111001: pixel[2:0] = 3'b000;
      14'b10011101111010: pixel[2:0] = 3'b000;
      14'b10011101111011: pixel[2:0] = 3'b000;
      14'b10011101111100: pixel[2:0] = 3'b000;
      14'b10011101111101: pixel[2:0] = 3'b000;
      14'b10011101111110: pixel[2:0] = 3'b111;
      14'b10011101111111: pixel[2:0] = 3'b111;
      14'b10011110000000: pixel[2:0] = 3'b111;
      14'b10011110000001: pixel[2:0] = 3'b111;
      14'b10011110000010: pixel[2:0] = 3'b111;
      14'b10011110000011: pixel[2:0] = 3'b000;
      14'b10011110000100: pixel[2:0] = 3'b000;
      14'b10011110000101: pixel[2:0] = 3'b000;
      14'b10011110000110: pixel[2:0] = 3'b000;
      14'b10011110000111: pixel[2:0] = 3'b000;
      14'b10100000000000: pixel[2:0] = 3'b000;
      14'b10100000000001: pixel[2:0] = 3'b000;
      14'b10100000000010: pixel[2:0] = 3'b111;
      14'b10100000000011: pixel[2:0] = 3'b111;
      14'b10100000000100: pixel[2:0] = 3'b111;
      14'b10100000000101: pixel[2:0] = 3'b111;
      14'b10100000000110: pixel[2:0] = 3'b111;
      14'b10100000000111: pixel[2:0] = 3'b000;
      14'b10100000001000: pixel[2:0] = 3'b000;
      14'b10100000001001: pixel[2:0] = 3'b000;
      14'b10100000001010: pixel[2:0] = 3'b000;
      14'b10100000001011: pixel[2:0] = 3'b000;
      14'b10100000001100: pixel[2:0] = 3'b000;
      14'b10100000001101: pixel[2:0] = 3'b000;
      14'b10100000001110: pixel[2:0] = 3'b000;
      14'b10100000001111: pixel[2:0] = 3'b000;
      14'b10100000010000: pixel[2:0] = 3'b000;
      14'b10100000010001: pixel[2:0] = 3'b000;
      14'b10100000010010: pixel[2:0] = 3'b000;
      14'b10100000010011: pixel[2:0] = 3'b000;
      14'b10100000010100: pixel[2:0] = 3'b000;
      14'b10100000010101: pixel[2:0] = 3'b000;
      14'b10100000010110: pixel[2:0] = 3'b000;
      14'b10100000010111: pixel[2:0] = 3'b000;
      14'b10100000011000: pixel[2:0] = 3'b000;
      14'b10100000011001: pixel[2:0] = 3'b111;
      14'b10100000011010: pixel[2:0] = 3'b111;
      14'b10100000011011: pixel[2:0] = 3'b111;
      14'b10100000011100: pixel[2:0] = 3'b111;
      14'b10100000011101: pixel[2:0] = 3'b111;
      14'b10100000011110: pixel[2:0] = 3'b111;
      14'b10100000011111: pixel[2:0] = 3'b111;
      14'b10100000100000: pixel[2:0] = 3'b111;
      14'b10100000100001: pixel[2:0] = 3'b111;
      14'b10100000100010: pixel[2:0] = 3'b111;
      14'b10100000100011: pixel[2:0] = 3'b111;
      14'b10100000100100: pixel[2:0] = 3'b111;
      14'b10100000100101: pixel[2:0] = 3'b111;
      14'b10100000100110: pixel[2:0] = 3'b111;
      14'b10100000100111: pixel[2:0] = 3'b111;
      14'b10100000101000: pixel[2:0] = 3'b111;
      14'b10100000101001: pixel[2:0] = 3'b111;
      14'b10100000101010: pixel[2:0] = 3'b000;
      14'b10100000101011: pixel[2:0] = 3'b000;
      14'b10100000101100: pixel[2:0] = 3'b000;
      14'b10100000101101: pixel[2:0] = 3'b111;
      14'b10100000101110: pixel[2:0] = 3'b111;
      14'b10100000101111: pixel[2:0] = 3'b111;
      14'b10100000110000: pixel[2:0] = 3'b111;
      14'b10100000110001: pixel[2:0] = 3'b111;
      14'b10100000110010: pixel[2:0] = 3'b000;
      14'b10100000110011: pixel[2:0] = 3'b000;
      14'b10100000110100: pixel[2:0] = 3'b000;
      14'b10100000110101: pixel[2:0] = 3'b000;
      14'b10100000110110: pixel[2:0] = 3'b000;
      14'b10100000110111: pixel[2:0] = 3'b000;
      14'b10100000111000: pixel[2:0] = 3'b000;
      14'b10100000111001: pixel[2:0] = 3'b000;
      14'b10100000111010: pixel[2:0] = 3'b000;
      14'b10100000111011: pixel[2:0] = 3'b000;
      14'b10100000111100: pixel[2:0] = 3'b000;
      14'b10100000111101: pixel[2:0] = 3'b000;
      14'b10100000111110: pixel[2:0] = 3'b111;
      14'b10100000111111: pixel[2:0] = 3'b111;
      14'b10100001000000: pixel[2:0] = 3'b111;
      14'b10100001000001: pixel[2:0] = 3'b111;
      14'b10100001000010: pixel[2:0] = 3'b000;
      14'b10100001000011: pixel[2:0] = 3'b000;
      14'b10100001000100: pixel[2:0] = 3'b000;
      14'b10100001000101: pixel[2:0] = 3'b000;
      14'b10100001000110: pixel[2:0] = 3'b000;
      14'b10100001000111: pixel[2:0] = 3'b000;
      14'b10100001001000: pixel[2:0] = 3'b000;
      14'b10100001001001: pixel[2:0] = 3'b111;
      14'b10100001001010: pixel[2:0] = 3'b111;
      14'b10100001001011: pixel[2:0] = 3'b111;
      14'b10100001001100: pixel[2:0] = 3'b111;
      14'b10100001001101: pixel[2:0] = 3'b111;
      14'b10100001001110: pixel[2:0] = 3'b000;
      14'b10100001001111: pixel[2:0] = 3'b000;
      14'b10100001010000: pixel[2:0] = 3'b000;
      14'b10100001010001: pixel[2:0] = 3'b000;
      14'b10100001010010: pixel[2:0] = 3'b000;
      14'b10100001010011: pixel[2:0] = 3'b000;
      14'b10100001010100: pixel[2:0] = 3'b000;
      14'b10100001010101: pixel[2:0] = 3'b000;
      14'b10100001010110: pixel[2:0] = 3'b000;
      14'b10100001010111: pixel[2:0] = 3'b000;
      14'b10100001011000: pixel[2:0] = 3'b000;
      14'b10100001011001: pixel[2:0] = 3'b000;
      14'b10100001011010: pixel[2:0] = 3'b111;
      14'b10100001011011: pixel[2:0] = 3'b111;
      14'b10100001011100: pixel[2:0] = 3'b111;
      14'b10100001011101: pixel[2:0] = 3'b111;
      14'b10100001011110: pixel[2:0] = 3'b111;
      14'b10100001011111: pixel[2:0] = 3'b111;
      14'b10100001100000: pixel[2:0] = 3'b111;
      14'b10100001100001: pixel[2:0] = 3'b111;
      14'b10100001100010: pixel[2:0] = 3'b111;
      14'b10100001100011: pixel[2:0] = 3'b111;
      14'b10100001100100: pixel[2:0] = 3'b111;
      14'b10100001100101: pixel[2:0] = 3'b111;
      14'b10100001100110: pixel[2:0] = 3'b111;
      14'b10100001100111: pixel[2:0] = 3'b111;
      14'b10100001101000: pixel[2:0] = 3'b111;
      14'b10100001101001: pixel[2:0] = 3'b111;
      14'b10100001101010: pixel[2:0] = 3'b111;
      14'b10100001101011: pixel[2:0] = 3'b000;
      14'b10100001101100: pixel[2:0] = 3'b000;
      14'b10100001101101: pixel[2:0] = 3'b000;
      14'b10100001101110: pixel[2:0] = 3'b000;
      14'b10100001101111: pixel[2:0] = 3'b000;
      14'b10100001110000: pixel[2:0] = 3'b111;
      14'b10100001110001: pixel[2:0] = 3'b111;
      14'b10100001110010: pixel[2:0] = 3'b111;
      14'b10100001110011: pixel[2:0] = 3'b111;
      14'b10100001110100: pixel[2:0] = 3'b111;
      14'b10100001110101: pixel[2:0] = 3'b000;
      14'b10100001110110: pixel[2:0] = 3'b000;
      14'b10100001110111: pixel[2:0] = 3'b000;
      14'b10100001111000: pixel[2:0] = 3'b000;
      14'b10100001111001: pixel[2:0] = 3'b000;
      14'b10100001111010: pixel[2:0] = 3'b000;
      14'b10100001111011: pixel[2:0] = 3'b000;
      14'b10100001111100: pixel[2:0] = 3'b000;
      14'b10100001111101: pixel[2:0] = 3'b000;
      14'b10100001111110: pixel[2:0] = 3'b111;
      14'b10100001111111: pixel[2:0] = 3'b111;
      14'b10100010000000: pixel[2:0] = 3'b111;
      14'b10100010000001: pixel[2:0] = 3'b111;
      14'b10100010000010: pixel[2:0] = 3'b111;
      14'b10100010000011: pixel[2:0] = 3'b111;
      14'b10100010000100: pixel[2:0] = 3'b000;
      14'b10100010000101: pixel[2:0] = 3'b000;
      14'b10100010000110: pixel[2:0] = 3'b000;
      14'b10100010000111: pixel[2:0] = 3'b000;
      14'b10100100000000: pixel[2:0] = 3'b000;
      14'b10100100000001: pixel[2:0] = 3'b000;
      14'b10100100000010: pixel[2:0] = 3'b111;
      14'b10100100000011: pixel[2:0] = 3'b111;
      14'b10100100000100: pixel[2:0] = 3'b111;
      14'b10100100000101: pixel[2:0] = 3'b111;
      14'b10100100000110: pixel[2:0] = 3'b111;
      14'b10100100000111: pixel[2:0] = 3'b000;
      14'b10100100001000: pixel[2:0] = 3'b000;
      14'b10100100001001: pixel[2:0] = 3'b000;
      14'b10100100001010: pixel[2:0] = 3'b000;
      14'b10100100001011: pixel[2:0] = 3'b000;
      14'b10100100001100: pixel[2:0] = 3'b000;
      14'b10100100001101: pixel[2:0] = 3'b000;
      14'b10100100001110: pixel[2:0] = 3'b000;
      14'b10100100001111: pixel[2:0] = 3'b000;
      14'b10100100010000: pixel[2:0] = 3'b000;
      14'b10100100010001: pixel[2:0] = 3'b000;
      14'b10100100010010: pixel[2:0] = 3'b000;
      14'b10100100010011: pixel[2:0] = 3'b000;
      14'b10100100010100: pixel[2:0] = 3'b000;
      14'b10100100010101: pixel[2:0] = 3'b000;
      14'b10100100010110: pixel[2:0] = 3'b000;
      14'b10100100010111: pixel[2:0] = 3'b000;
      14'b10100100011000: pixel[2:0] = 3'b000;
      14'b10100100011001: pixel[2:0] = 3'b111;
      14'b10100100011010: pixel[2:0] = 3'b111;
      14'b10100100011011: pixel[2:0] = 3'b111;
      14'b10100100011100: pixel[2:0] = 3'b111;
      14'b10100100011101: pixel[2:0] = 3'b111;
      14'b10100100011110: pixel[2:0] = 3'b111;
      14'b10100100011111: pixel[2:0] = 3'b111;
      14'b10100100100000: pixel[2:0] = 3'b111;
      14'b10100100100001: pixel[2:0] = 3'b111;
      14'b10100100100010: pixel[2:0] = 3'b111;
      14'b10100100100011: pixel[2:0] = 3'b111;
      14'b10100100100100: pixel[2:0] = 3'b111;
      14'b10100100100101: pixel[2:0] = 3'b111;
      14'b10100100100110: pixel[2:0] = 3'b111;
      14'b10100100100111: pixel[2:0] = 3'b111;
      14'b10100100101000: pixel[2:0] = 3'b111;
      14'b10100100101001: pixel[2:0] = 3'b111;
      14'b10100100101010: pixel[2:0] = 3'b000;
      14'b10100100101011: pixel[2:0] = 3'b000;
      14'b10100100101100: pixel[2:0] = 3'b000;
      14'b10100100101101: pixel[2:0] = 3'b111;
      14'b10100100101110: pixel[2:0] = 3'b111;
      14'b10100100101111: pixel[2:0] = 3'b111;
      14'b10100100110000: pixel[2:0] = 3'b111;
      14'b10100100110001: pixel[2:0] = 3'b111;
      14'b10100100110010: pixel[2:0] = 3'b000;
      14'b10100100110011: pixel[2:0] = 3'b000;
      14'b10100100110100: pixel[2:0] = 3'b000;
      14'b10100100110101: pixel[2:0] = 3'b000;
      14'b10100100110110: pixel[2:0] = 3'b000;
      14'b10100100110111: pixel[2:0] = 3'b000;
      14'b10100100111000: pixel[2:0] = 3'b000;
      14'b10100100111001: pixel[2:0] = 3'b000;
      14'b10100100111010: pixel[2:0] = 3'b000;
      14'b10100100111011: pixel[2:0] = 3'b000;
      14'b10100100111100: pixel[2:0] = 3'b000;
      14'b10100100111101: pixel[2:0] = 3'b000;
      14'b10100100111110: pixel[2:0] = 3'b111;
      14'b10100100111111: pixel[2:0] = 3'b111;
      14'b10100101000000: pixel[2:0] = 3'b111;
      14'b10100101000001: pixel[2:0] = 3'b111;
      14'b10100101000010: pixel[2:0] = 3'b111;
      14'b10100101000011: pixel[2:0] = 3'b000;
      14'b10100101000100: pixel[2:0] = 3'b000;
      14'b10100101000101: pixel[2:0] = 3'b000;
      14'b10100101000110: pixel[2:0] = 3'b000;
      14'b10100101000111: pixel[2:0] = 3'b000;
      14'b10100101001000: pixel[2:0] = 3'b000;
      14'b10100101001001: pixel[2:0] = 3'b111;
      14'b10100101001010: pixel[2:0] = 3'b111;
      14'b10100101001011: pixel[2:0] = 3'b111;
      14'b10100101001100: pixel[2:0] = 3'b111;
      14'b10100101001101: pixel[2:0] = 3'b111;
      14'b10100101001110: pixel[2:0] = 3'b000;
      14'b10100101001111: pixel[2:0] = 3'b000;
      14'b10100101010000: pixel[2:0] = 3'b000;
      14'b10100101010001: pixel[2:0] = 3'b000;
      14'b10100101010010: pixel[2:0] = 3'b000;
      14'b10100101010011: pixel[2:0] = 3'b000;
      14'b10100101010100: pixel[2:0] = 3'b000;
      14'b10100101010101: pixel[2:0] = 3'b000;
      14'b10100101010110: pixel[2:0] = 3'b000;
      14'b10100101010111: pixel[2:0] = 3'b000;
      14'b10100101011000: pixel[2:0] = 3'b000;
      14'b10100101011001: pixel[2:0] = 3'b000;
      14'b10100101011010: pixel[2:0] = 3'b111;
      14'b10100101011011: pixel[2:0] = 3'b111;
      14'b10100101011100: pixel[2:0] = 3'b111;
      14'b10100101011101: pixel[2:0] = 3'b111;
      14'b10100101011110: pixel[2:0] = 3'b111;
      14'b10100101011111: pixel[2:0] = 3'b111;
      14'b10100101100000: pixel[2:0] = 3'b111;
      14'b10100101100001: pixel[2:0] = 3'b111;
      14'b10100101100010: pixel[2:0] = 3'b111;
      14'b10100101100011: pixel[2:0] = 3'b111;
      14'b10100101100100: pixel[2:0] = 3'b111;
      14'b10100101100101: pixel[2:0] = 3'b111;
      14'b10100101100110: pixel[2:0] = 3'b111;
      14'b10100101100111: pixel[2:0] = 3'b111;
      14'b10100101101000: pixel[2:0] = 3'b111;
      14'b10100101101001: pixel[2:0] = 3'b111;
      14'b10100101101010: pixel[2:0] = 3'b111;
      14'b10100101101011: pixel[2:0] = 3'b000;
      14'b10100101101100: pixel[2:0] = 3'b000;
      14'b10100101101101: pixel[2:0] = 3'b000;
      14'b10100101101110: pixel[2:0] = 3'b000;
      14'b10100101101111: pixel[2:0] = 3'b000;
      14'b10100101110000: pixel[2:0] = 3'b111;
      14'b10100101110001: pixel[2:0] = 3'b111;
      14'b10100101110010: pixel[2:0] = 3'b111;
      14'b10100101110011: pixel[2:0] = 3'b111;
      14'b10100101110100: pixel[2:0] = 3'b111;
      14'b10100101110101: pixel[2:0] = 3'b000;
      14'b10100101110110: pixel[2:0] = 3'b000;
      14'b10100101110111: pixel[2:0] = 3'b000;
      14'b10100101111000: pixel[2:0] = 3'b000;
      14'b10100101111001: pixel[2:0] = 3'b000;
      14'b10100101111010: pixel[2:0] = 3'b000;
      14'b10100101111011: pixel[2:0] = 3'b000;
      14'b10100101111100: pixel[2:0] = 3'b000;
      14'b10100101111101: pixel[2:0] = 3'b000;
      14'b10100101111110: pixel[2:0] = 3'b000;
      14'b10100101111111: pixel[2:0] = 3'b111;
      14'b10100110000000: pixel[2:0] = 3'b111;
      14'b10100110000001: pixel[2:0] = 3'b111;
      14'b10100110000010: pixel[2:0] = 3'b111;
      14'b10100110000011: pixel[2:0] = 3'b111;
      14'b10100110000100: pixel[2:0] = 3'b000;
      14'b10100110000101: pixel[2:0] = 3'b000;
      14'b10100110000110: pixel[2:0] = 3'b000;
      14'b10100110000111: pixel[2:0] = 3'b000;
      14'b10101000000000: pixel[2:0] = 3'b000;
      14'b10101000000001: pixel[2:0] = 3'b000;
      14'b10101000000010: pixel[2:0] = 3'b111;
      14'b10101000000011: pixel[2:0] = 3'b111;
      14'b10101000000100: pixel[2:0] = 3'b111;
      14'b10101000000101: pixel[2:0] = 3'b111;
      14'b10101000000110: pixel[2:0] = 3'b111;
      14'b10101000000111: pixel[2:0] = 3'b000;
      14'b10101000001000: pixel[2:0] = 3'b000;
      14'b10101000001001: pixel[2:0] = 3'b000;
      14'b10101000001010: pixel[2:0] = 3'b000;
      14'b10101000001011: pixel[2:0] = 3'b000;
      14'b10101000001100: pixel[2:0] = 3'b000;
      14'b10101000001101: pixel[2:0] = 3'b000;
      14'b10101000001110: pixel[2:0] = 3'b000;
      14'b10101000001111: pixel[2:0] = 3'b000;
      14'b10101000010000: pixel[2:0] = 3'b000;
      14'b10101000010001: pixel[2:0] = 3'b000;
      14'b10101000010010: pixel[2:0] = 3'b000;
      14'b10101000010011: pixel[2:0] = 3'b000;
      14'b10101000010100: pixel[2:0] = 3'b000;
      14'b10101000010101: pixel[2:0] = 3'b000;
      14'b10101000010110: pixel[2:0] = 3'b000;
      14'b10101000010111: pixel[2:0] = 3'b000;
      14'b10101000011000: pixel[2:0] = 3'b000;
      14'b10101000011001: pixel[2:0] = 3'b111;
      14'b10101000011010: pixel[2:0] = 3'b111;
      14'b10101000011011: pixel[2:0] = 3'b111;
      14'b10101000011100: pixel[2:0] = 3'b111;
      14'b10101000011101: pixel[2:0] = 3'b111;
      14'b10101000011110: pixel[2:0] = 3'b111;
      14'b10101000011111: pixel[2:0] = 3'b111;
      14'b10101000100000: pixel[2:0] = 3'b111;
      14'b10101000100001: pixel[2:0] = 3'b111;
      14'b10101000100010: pixel[2:0] = 3'b111;
      14'b10101000100011: pixel[2:0] = 3'b111;
      14'b10101000100100: pixel[2:0] = 3'b111;
      14'b10101000100101: pixel[2:0] = 3'b111;
      14'b10101000100110: pixel[2:0] = 3'b111;
      14'b10101000100111: pixel[2:0] = 3'b111;
      14'b10101000101000: pixel[2:0] = 3'b111;
      14'b10101000101001: pixel[2:0] = 3'b111;
      14'b10101000101010: pixel[2:0] = 3'b000;
      14'b10101000101011: pixel[2:0] = 3'b000;
      14'b10101000101100: pixel[2:0] = 3'b000;
      14'b10101000101101: pixel[2:0] = 3'b111;
      14'b10101000101110: pixel[2:0] = 3'b111;
      14'b10101000101111: pixel[2:0] = 3'b111;
      14'b10101000110000: pixel[2:0] = 3'b111;
      14'b10101000110001: pixel[2:0] = 3'b111;
      14'b10101000110010: pixel[2:0] = 3'b000;
      14'b10101000110011: pixel[2:0] = 3'b000;
      14'b10101000110100: pixel[2:0] = 3'b000;
      14'b10101000110101: pixel[2:0] = 3'b000;
      14'b10101000110110: pixel[2:0] = 3'b000;
      14'b10101000110111: pixel[2:0] = 3'b000;
      14'b10101000111000: pixel[2:0] = 3'b000;
      14'b10101000111001: pixel[2:0] = 3'b000;
      14'b10101000111010: pixel[2:0] = 3'b000;
      14'b10101000111011: pixel[2:0] = 3'b000;
      14'b10101000111100: pixel[2:0] = 3'b000;
      14'b10101000111101: pixel[2:0] = 3'b000;
      14'b10101000111110: pixel[2:0] = 3'b111;
      14'b10101000111111: pixel[2:0] = 3'b111;
      14'b10101001000000: pixel[2:0] = 3'b111;
      14'b10101001000001: pixel[2:0] = 3'b111;
      14'b10101001000010: pixel[2:0] = 3'b111;
      14'b10101001000011: pixel[2:0] = 3'b000;
      14'b10101001000100: pixel[2:0] = 3'b000;
      14'b10101001000101: pixel[2:0] = 3'b000;
      14'b10101001000110: pixel[2:0] = 3'b000;
      14'b10101001000111: pixel[2:0] = 3'b000;
      14'b10101001001000: pixel[2:0] = 3'b000;
      14'b10101001001001: pixel[2:0] = 3'b111;
      14'b10101001001010: pixel[2:0] = 3'b111;
      14'b10101001001011: pixel[2:0] = 3'b111;
      14'b10101001001100: pixel[2:0] = 3'b111;
      14'b10101001001101: pixel[2:0] = 3'b111;
      14'b10101001001110: pixel[2:0] = 3'b000;
      14'b10101001001111: pixel[2:0] = 3'b000;
      14'b10101001010000: pixel[2:0] = 3'b000;
      14'b10101001010001: pixel[2:0] = 3'b000;
      14'b10101001010010: pixel[2:0] = 3'b000;
      14'b10101001010011: pixel[2:0] = 3'b000;
      14'b10101001010100: pixel[2:0] = 3'b000;
      14'b10101001010101: pixel[2:0] = 3'b000;
      14'b10101001010110: pixel[2:0] = 3'b000;
      14'b10101001010111: pixel[2:0] = 3'b000;
      14'b10101001011000: pixel[2:0] = 3'b000;
      14'b10101001011001: pixel[2:0] = 3'b000;
      14'b10101001011010: pixel[2:0] = 3'b111;
      14'b10101001011011: pixel[2:0] = 3'b111;
      14'b10101001011100: pixel[2:0] = 3'b111;
      14'b10101001011101: pixel[2:0] = 3'b111;
      14'b10101001011110: pixel[2:0] = 3'b111;
      14'b10101001011111: pixel[2:0] = 3'b111;
      14'b10101001100000: pixel[2:0] = 3'b111;
      14'b10101001100001: pixel[2:0] = 3'b111;
      14'b10101001100010: pixel[2:0] = 3'b111;
      14'b10101001100011: pixel[2:0] = 3'b111;
      14'b10101001100100: pixel[2:0] = 3'b111;
      14'b10101001100101: pixel[2:0] = 3'b111;
      14'b10101001100110: pixel[2:0] = 3'b111;
      14'b10101001100111: pixel[2:0] = 3'b111;
      14'b10101001101000: pixel[2:0] = 3'b111;
      14'b10101001101001: pixel[2:0] = 3'b111;
      14'b10101001101010: pixel[2:0] = 3'b111;
      14'b10101001101011: pixel[2:0] = 3'b000;
      14'b10101001101100: pixel[2:0] = 3'b000;
      14'b10101001101101: pixel[2:0] = 3'b000;
      14'b10101001101110: pixel[2:0] = 3'b000;
      14'b10101001101111: pixel[2:0] = 3'b000;
      14'b10101001110000: pixel[2:0] = 3'b111;
      14'b10101001110001: pixel[2:0] = 3'b111;
      14'b10101001110010: pixel[2:0] = 3'b111;
      14'b10101001110011: pixel[2:0] = 3'b111;
      14'b10101001110100: pixel[2:0] = 3'b111;
      14'b10101001110101: pixel[2:0] = 3'b000;
      14'b10101001110110: pixel[2:0] = 3'b000;
      14'b10101001110111: pixel[2:0] = 3'b000;
      14'b10101001111000: pixel[2:0] = 3'b000;
      14'b10101001111001: pixel[2:0] = 3'b000;
      14'b10101001111010: pixel[2:0] = 3'b000;
      14'b10101001111011: pixel[2:0] = 3'b000;
      14'b10101001111100: pixel[2:0] = 3'b000;
      14'b10101001111101: pixel[2:0] = 3'b000;
      14'b10101001111110: pixel[2:0] = 3'b000;
      14'b10101001111111: pixel[2:0] = 3'b111;
      14'b10101010000000: pixel[2:0] = 3'b111;
      14'b10101010000001: pixel[2:0] = 3'b111;
      14'b10101010000010: pixel[2:0] = 3'b111;
      14'b10101010000011: pixel[2:0] = 3'b111;
      14'b10101010000100: pixel[2:0] = 3'b000;
      14'b10101010000101: pixel[2:0] = 3'b000;
      14'b10101010000110: pixel[2:0] = 3'b000;
      14'b10101010000111: pixel[2:0] = 3'b000;
      14'b10101100000000: pixel[2:0] = 3'b000;
      14'b10101100000001: pixel[2:0] = 3'b000;
      14'b10101100000010: pixel[2:0] = 3'b000;
      14'b10101100000011: pixel[2:0] = 3'b000;
      14'b10101100000100: pixel[2:0] = 3'b000;
      14'b10101100000101: pixel[2:0] = 3'b000;
      14'b10101100000110: pixel[2:0] = 3'b000;
      14'b10101100000111: pixel[2:0] = 3'b000;
      14'b10101100001000: pixel[2:0] = 3'b000;
      14'b10101100001001: pixel[2:0] = 3'b000;
      14'b10101100001010: pixel[2:0] = 3'b000;
      14'b10101100001011: pixel[2:0] = 3'b000;
      14'b10101100001100: pixel[2:0] = 3'b000;
      14'b10101100001101: pixel[2:0] = 3'b000;
      14'b10101100001110: pixel[2:0] = 3'b000;
      14'b10101100001111: pixel[2:0] = 3'b000;
      14'b10101100010000: pixel[2:0] = 3'b000;
      14'b10101100010001: pixel[2:0] = 3'b000;
      14'b10101100010010: pixel[2:0] = 3'b000;
      14'b10101100010011: pixel[2:0] = 3'b000;
      14'b10101100010100: pixel[2:0] = 3'b000;
      14'b10101100010101: pixel[2:0] = 3'b000;
      14'b10101100010110: pixel[2:0] = 3'b000;
      14'b10101100010111: pixel[2:0] = 3'b000;
      14'b10101100011000: pixel[2:0] = 3'b000;
      14'b10101100011001: pixel[2:0] = 3'b000;
      14'b10101100011010: pixel[2:0] = 3'b000;
      14'b10101100011011: pixel[2:0] = 3'b000;
      14'b10101100011100: pixel[2:0] = 3'b000;
      14'b10101100011101: pixel[2:0] = 3'b000;
      14'b10101100011110: pixel[2:0] = 3'b000;
      14'b10101100011111: pixel[2:0] = 3'b000;
      14'b10101100100000: pixel[2:0] = 3'b000;
      14'b10101100100001: pixel[2:0] = 3'b000;
      14'b10101100100010: pixel[2:0] = 3'b000;
      14'b10101100100011: pixel[2:0] = 3'b000;
      14'b10101100100100: pixel[2:0] = 3'b000;
      14'b10101100100101: pixel[2:0] = 3'b000;
      14'b10101100100110: pixel[2:0] = 3'b000;
      14'b10101100100111: pixel[2:0] = 3'b000;
      14'b10101100101000: pixel[2:0] = 3'b000;
      14'b10101100101001: pixel[2:0] = 3'b000;
      14'b10101100101010: pixel[2:0] = 3'b000;
      14'b10101100101011: pixel[2:0] = 3'b000;
      14'b10101100101100: pixel[2:0] = 3'b000;
      14'b10101100101101: pixel[2:0] = 3'b000;
      14'b10101100101110: pixel[2:0] = 3'b000;
      14'b10101100101111: pixel[2:0] = 3'b000;
      14'b10101100110000: pixel[2:0] = 3'b000;
      14'b10101100110001: pixel[2:0] = 3'b000;
      14'b10101100110010: pixel[2:0] = 3'b000;
      14'b10101100110011: pixel[2:0] = 3'b000;
      14'b10101100110100: pixel[2:0] = 3'b000;
      14'b10101100110101: pixel[2:0] = 3'b000;
      14'b10101100110110: pixel[2:0] = 3'b000;
      14'b10101100110111: pixel[2:0] = 3'b000;
      14'b10101100111000: pixel[2:0] = 3'b000;
      14'b10101100111001: pixel[2:0] = 3'b000;
      14'b10101100111010: pixel[2:0] = 3'b000;
      14'b10101100111011: pixel[2:0] = 3'b000;
      14'b10101100111100: pixel[2:0] = 3'b000;
      14'b10101100111101: pixel[2:0] = 3'b000;
      14'b10101100111110: pixel[2:0] = 3'b000;
      14'b10101100111111: pixel[2:0] = 3'b000;
      14'b10101101000000: pixel[2:0] = 3'b000;
      14'b10101101000001: pixel[2:0] = 3'b000;
      14'b10101101000010: pixel[2:0] = 3'b000;
      14'b10101101000011: pixel[2:0] = 3'b000;
      14'b10101101000100: pixel[2:0] = 3'b000;
      14'b10101101000101: pixel[2:0] = 3'b000;
      14'b10101101000110: pixel[2:0] = 3'b000;
      14'b10101101000111: pixel[2:0] = 3'b000;
      14'b10101101001000: pixel[2:0] = 3'b000;
      14'b10101101001001: pixel[2:0] = 3'b000;
      14'b10101101001010: pixel[2:0] = 3'b000;
      14'b10101101001011: pixel[2:0] = 3'b000;
      14'b10101101001100: pixel[2:0] = 3'b000;
      14'b10101101001101: pixel[2:0] = 3'b000;
      14'b10101101001110: pixel[2:0] = 3'b000;
      14'b10101101001111: pixel[2:0] = 3'b000;
      14'b10101101010000: pixel[2:0] = 3'b000;
      14'b10101101010001: pixel[2:0] = 3'b000;
      14'b10101101010010: pixel[2:0] = 3'b000;
      14'b10101101010011: pixel[2:0] = 3'b000;
      14'b10101101010100: pixel[2:0] = 3'b000;
      14'b10101101010101: pixel[2:0] = 3'b000;
      14'b10101101010110: pixel[2:0] = 3'b000;
      14'b10101101010111: pixel[2:0] = 3'b000;
      14'b10101101011000: pixel[2:0] = 3'b000;
      14'b10101101011001: pixel[2:0] = 3'b000;
      14'b10101101011010: pixel[2:0] = 3'b000;
      14'b10101101011011: pixel[2:0] = 3'b000;
      14'b10101101011100: pixel[2:0] = 3'b000;
      14'b10101101011101: pixel[2:0] = 3'b000;
      14'b10101101011110: pixel[2:0] = 3'b000;
      14'b10101101011111: pixel[2:0] = 3'b000;
      14'b10101101100000: pixel[2:0] = 3'b000;
      14'b10101101100001: pixel[2:0] = 3'b000;
      14'b10101101100010: pixel[2:0] = 3'b000;
      14'b10101101100011: pixel[2:0] = 3'b000;
      14'b10101101100100: pixel[2:0] = 3'b000;
      14'b10101101100101: pixel[2:0] = 3'b000;
      14'b10101101100110: pixel[2:0] = 3'b000;
      14'b10101101100111: pixel[2:0] = 3'b000;
      14'b10101101101000: pixel[2:0] = 3'b000;
      14'b10101101101001: pixel[2:0] = 3'b000;
      14'b10101101101010: pixel[2:0] = 3'b000;
      14'b10101101101011: pixel[2:0] = 3'b000;
      14'b10101101101100: pixel[2:0] = 3'b000;
      14'b10101101101101: pixel[2:0] = 3'b000;
      14'b10101101101110: pixel[2:0] = 3'b000;
      14'b10101101101111: pixel[2:0] = 3'b000;
      14'b10101101110000: pixel[2:0] = 3'b000;
      14'b10101101110001: pixel[2:0] = 3'b000;
      14'b10101101110010: pixel[2:0] = 3'b000;
      14'b10101101110011: pixel[2:0] = 3'b000;
      14'b10101101110100: pixel[2:0] = 3'b000;
      14'b10101101110101: pixel[2:0] = 3'b000;
      14'b10101101110110: pixel[2:0] = 3'b000;
      14'b10101101110111: pixel[2:0] = 3'b000;
      14'b10101101111000: pixel[2:0] = 3'b000;
      14'b10101101111001: pixel[2:0] = 3'b000;
      14'b10101101111010: pixel[2:0] = 3'b000;
      14'b10101101111011: pixel[2:0] = 3'b000;
      14'b10101101111100: pixel[2:0] = 3'b000;
      14'b10101101111101: pixel[2:0] = 3'b000;
      14'b10101101111110: pixel[2:0] = 3'b000;
      14'b10101101111111: pixel[2:0] = 3'b000;
      14'b10101110000000: pixel[2:0] = 3'b000;
      14'b10101110000001: pixel[2:0] = 3'b000;
      14'b10101110000010: pixel[2:0] = 3'b000;
      14'b10101110000011: pixel[2:0] = 3'b000;
      14'b10101110000100: pixel[2:0] = 3'b000;
      14'b10101110000101: pixel[2:0] = 3'b000;
      14'b10101110000110: pixel[2:0] = 3'b000;
      14'b10101110000111: pixel[2:0] = 3'b000;
      14'b10110000000000: pixel[2:0] = 3'b000;
      14'b10110000000001: pixel[2:0] = 3'b000;
      14'b10110000000010: pixel[2:0] = 3'b000;
      14'b10110000000011: pixel[2:0] = 3'b000;
      14'b10110000000100: pixel[2:0] = 3'b000;
      14'b10110000000101: pixel[2:0] = 3'b000;
      14'b10110000000110: pixel[2:0] = 3'b000;
      14'b10110000000111: pixel[2:0] = 3'b000;
      14'b10110000001000: pixel[2:0] = 3'b000;
      14'b10110000001001: pixel[2:0] = 3'b000;
      14'b10110000001010: pixel[2:0] = 3'b000;
      14'b10110000001011: pixel[2:0] = 3'b000;
      14'b10110000001100: pixel[2:0] = 3'b000;
      14'b10110000001101: pixel[2:0] = 3'b000;
      14'b10110000001110: pixel[2:0] = 3'b000;
      14'b10110000001111: pixel[2:0] = 3'b000;
      14'b10110000010000: pixel[2:0] = 3'b000;
      14'b10110000010001: pixel[2:0] = 3'b000;
      14'b10110000010010: pixel[2:0] = 3'b000;
      14'b10110000010011: pixel[2:0] = 3'b000;
      14'b10110000010100: pixel[2:0] = 3'b000;
      14'b10110000010101: pixel[2:0] = 3'b000;
      14'b10110000010110: pixel[2:0] = 3'b000;
      14'b10110000010111: pixel[2:0] = 3'b000;
      14'b10110000011000: pixel[2:0] = 3'b000;
      14'b10110000011001: pixel[2:0] = 3'b000;
      14'b10110000011010: pixel[2:0] = 3'b000;
      14'b10110000011011: pixel[2:0] = 3'b000;
      14'b10110000011100: pixel[2:0] = 3'b000;
      14'b10110000011101: pixel[2:0] = 3'b000;
      14'b10110000011110: pixel[2:0] = 3'b000;
      14'b10110000011111: pixel[2:0] = 3'b000;
      14'b10110000100000: pixel[2:0] = 3'b000;
      14'b10110000100001: pixel[2:0] = 3'b000;
      14'b10110000100010: pixel[2:0] = 3'b000;
      14'b10110000100011: pixel[2:0] = 3'b000;
      14'b10110000100100: pixel[2:0] = 3'b000;
      14'b10110000100101: pixel[2:0] = 3'b000;
      14'b10110000100110: pixel[2:0] = 3'b000;
      14'b10110000100111: pixel[2:0] = 3'b000;
      14'b10110000101000: pixel[2:0] = 3'b000;
      14'b10110000101001: pixel[2:0] = 3'b000;
      14'b10110000101010: pixel[2:0] = 3'b000;
      14'b10110000101011: pixel[2:0] = 3'b000;
      14'b10110000101100: pixel[2:0] = 3'b000;
      14'b10110000101101: pixel[2:0] = 3'b000;
      14'b10110000101110: pixel[2:0] = 3'b000;
      14'b10110000101111: pixel[2:0] = 3'b000;
      14'b10110000110000: pixel[2:0] = 3'b000;
      14'b10110000110001: pixel[2:0] = 3'b000;
      14'b10110000110010: pixel[2:0] = 3'b000;
      14'b10110000110011: pixel[2:0] = 3'b000;
      14'b10110000110100: pixel[2:0] = 3'b000;
      14'b10110000110101: pixel[2:0] = 3'b000;
      14'b10110000110110: pixel[2:0] = 3'b000;
      14'b10110000110111: pixel[2:0] = 3'b000;
      14'b10110000111000: pixel[2:0] = 3'b000;
      14'b10110000111001: pixel[2:0] = 3'b000;
      14'b10110000111010: pixel[2:0] = 3'b000;
      14'b10110000111011: pixel[2:0] = 3'b000;
      14'b10110000111100: pixel[2:0] = 3'b000;
      14'b10110000111101: pixel[2:0] = 3'b000;
      14'b10110000111110: pixel[2:0] = 3'b000;
      14'b10110000111111: pixel[2:0] = 3'b000;
      14'b10110001000000: pixel[2:0] = 3'b000;
      14'b10110001000001: pixel[2:0] = 3'b000;
      14'b10110001000010: pixel[2:0] = 3'b000;
      14'b10110001000011: pixel[2:0] = 3'b000;
      14'b10110001000100: pixel[2:0] = 3'b000;
      14'b10110001000101: pixel[2:0] = 3'b000;
      14'b10110001000110: pixel[2:0] = 3'b000;
      14'b10110001000111: pixel[2:0] = 3'b000;
      14'b10110001001000: pixel[2:0] = 3'b000;
      14'b10110001001001: pixel[2:0] = 3'b000;
      14'b10110001001010: pixel[2:0] = 3'b000;
      14'b10110001001011: pixel[2:0] = 3'b000;
      14'b10110001001100: pixel[2:0] = 3'b000;
      14'b10110001001101: pixel[2:0] = 3'b000;
      14'b10110001001110: pixel[2:0] = 3'b000;
      14'b10110001001111: pixel[2:0] = 3'b000;
      14'b10110001010000: pixel[2:0] = 3'b000;
      14'b10110001010001: pixel[2:0] = 3'b000;
      14'b10110001010010: pixel[2:0] = 3'b000;
      14'b10110001010011: pixel[2:0] = 3'b000;
      14'b10110001010100: pixel[2:0] = 3'b000;
      14'b10110001010101: pixel[2:0] = 3'b000;
      14'b10110001010110: pixel[2:0] = 3'b000;
      14'b10110001010111: pixel[2:0] = 3'b000;
      14'b10110001011000: pixel[2:0] = 3'b000;
      14'b10110001011001: pixel[2:0] = 3'b000;
      14'b10110001011010: pixel[2:0] = 3'b000;
      14'b10110001011011: pixel[2:0] = 3'b000;
      14'b10110001011100: pixel[2:0] = 3'b000;
      14'b10110001011101: pixel[2:0] = 3'b000;
      14'b10110001011110: pixel[2:0] = 3'b000;
      14'b10110001011111: pixel[2:0] = 3'b000;
      14'b10110001100000: pixel[2:0] = 3'b000;
      14'b10110001100001: pixel[2:0] = 3'b000;
      14'b10110001100010: pixel[2:0] = 3'b000;
      14'b10110001100011: pixel[2:0] = 3'b000;
      14'b10110001100100: pixel[2:0] = 3'b000;
      14'b10110001100101: pixel[2:0] = 3'b000;
      14'b10110001100110: pixel[2:0] = 3'b000;
      14'b10110001100111: pixel[2:0] = 3'b000;
      14'b10110001101000: pixel[2:0] = 3'b000;
      14'b10110001101001: pixel[2:0] = 3'b000;
      14'b10110001101010: pixel[2:0] = 3'b000;
      14'b10110001101011: pixel[2:0] = 3'b000;
      14'b10110001101100: pixel[2:0] = 3'b000;
      14'b10110001101101: pixel[2:0] = 3'b000;
      14'b10110001101110: pixel[2:0] = 3'b000;
      14'b10110001101111: pixel[2:0] = 3'b000;
      14'b10110001110000: pixel[2:0] = 3'b000;
      14'b10110001110001: pixel[2:0] = 3'b000;
      14'b10110001110010: pixel[2:0] = 3'b000;
      14'b10110001110011: pixel[2:0] = 3'b000;
      14'b10110001110100: pixel[2:0] = 3'b000;
      14'b10110001110101: pixel[2:0] = 3'b000;
      14'b10110001110110: pixel[2:0] = 3'b000;
      14'b10110001110111: pixel[2:0] = 3'b000;
      14'b10110001111000: pixel[2:0] = 3'b000;
      14'b10110001111001: pixel[2:0] = 3'b000;
      14'b10110001111010: pixel[2:0] = 3'b000;
      14'b10110001111011: pixel[2:0] = 3'b000;
      14'b10110001111100: pixel[2:0] = 3'b000;
      14'b10110001111101: pixel[2:0] = 3'b000;
      14'b10110001111110: pixel[2:0] = 3'b000;
      14'b10110001111111: pixel[2:0] = 3'b000;
      14'b10110010000000: pixel[2:0] = 3'b000;
      14'b10110010000001: pixel[2:0] = 3'b000;
      14'b10110010000010: pixel[2:0] = 3'b000;
      14'b10110010000011: pixel[2:0] = 3'b000;
      14'b10110010000100: pixel[2:0] = 3'b000;
      14'b10110010000101: pixel[2:0] = 3'b000;
      14'b10110010000110: pixel[2:0] = 3'b000;
      14'b10110010000111: pixel[2:0] = 3'b000;
      14'b10110100000000: pixel[2:0] = 3'b000;
      14'b10110100000001: pixel[2:0] = 3'b000;
      14'b10110100000010: pixel[2:0] = 3'b000;
      14'b10110100000011: pixel[2:0] = 3'b000;
      14'b10110100000100: pixel[2:0] = 3'b000;
      14'b10110100000101: pixel[2:0] = 3'b000;
      14'b10110100000110: pixel[2:0] = 3'b000;
      14'b10110100000111: pixel[2:0] = 3'b000;
      14'b10110100001000: pixel[2:0] = 3'b000;
      14'b10110100001001: pixel[2:0] = 3'b000;
      14'b10110100001010: pixel[2:0] = 3'b000;
      14'b10110100001011: pixel[2:0] = 3'b000;
      14'b10110100001100: pixel[2:0] = 3'b000;
      14'b10110100001101: pixel[2:0] = 3'b000;
      14'b10110100001110: pixel[2:0] = 3'b000;
      14'b10110100001111: pixel[2:0] = 3'b000;
      14'b10110100010000: pixel[2:0] = 3'b000;
      14'b10110100010001: pixel[2:0] = 3'b000;
      14'b10110100010010: pixel[2:0] = 3'b000;
      14'b10110100010011: pixel[2:0] = 3'b000;
      14'b10110100010100: pixel[2:0] = 3'b000;
      14'b10110100010101: pixel[2:0] = 3'b000;
      14'b10110100010110: pixel[2:0] = 3'b000;
      14'b10110100010111: pixel[2:0] = 3'b000;
      14'b10110100011000: pixel[2:0] = 3'b000;
      14'b10110100011001: pixel[2:0] = 3'b000;
      14'b10110100011010: pixel[2:0] = 3'b000;
      14'b10110100011011: pixel[2:0] = 3'b000;
      14'b10110100011100: pixel[2:0] = 3'b000;
      14'b10110100011101: pixel[2:0] = 3'b000;
      14'b10110100011110: pixel[2:0] = 3'b000;
      14'b10110100011111: pixel[2:0] = 3'b000;
      14'b10110100100000: pixel[2:0] = 3'b000;
      14'b10110100100001: pixel[2:0] = 3'b000;
      14'b10110100100010: pixel[2:0] = 3'b000;
      14'b10110100100011: pixel[2:0] = 3'b000;
      14'b10110100100100: pixel[2:0] = 3'b000;
      14'b10110100100101: pixel[2:0] = 3'b000;
      14'b10110100100110: pixel[2:0] = 3'b000;
      14'b10110100100111: pixel[2:0] = 3'b000;
      14'b10110100101000: pixel[2:0] = 3'b000;
      14'b10110100101001: pixel[2:0] = 3'b000;
      14'b10110100101010: pixel[2:0] = 3'b000;
      14'b10110100101011: pixel[2:0] = 3'b000;
      14'b10110100101100: pixel[2:0] = 3'b000;
      14'b10110100101101: pixel[2:0] = 3'b000;
      14'b10110100101110: pixel[2:0] = 3'b000;
      14'b10110100101111: pixel[2:0] = 3'b000;
      14'b10110100110000: pixel[2:0] = 3'b000;
      14'b10110100110001: pixel[2:0] = 3'b000;
      14'b10110100110010: pixel[2:0] = 3'b000;
      14'b10110100110011: pixel[2:0] = 3'b000;
      14'b10110100110100: pixel[2:0] = 3'b000;
      14'b10110100110101: pixel[2:0] = 3'b000;
      14'b10110100110110: pixel[2:0] = 3'b000;
      14'b10110100110111: pixel[2:0] = 3'b000;
      14'b10110100111000: pixel[2:0] = 3'b000;
      14'b10110100111001: pixel[2:0] = 3'b000;
      14'b10110100111010: pixel[2:0] = 3'b000;
      14'b10110100111011: pixel[2:0] = 3'b000;
      14'b10110100111100: pixel[2:0] = 3'b000;
      14'b10110100111101: pixel[2:0] = 3'b000;
      14'b10110100111110: pixel[2:0] = 3'b000;
      14'b10110100111111: pixel[2:0] = 3'b000;
      14'b10110101000000: pixel[2:0] = 3'b000;
      14'b10110101000001: pixel[2:0] = 3'b000;
      14'b10110101000010: pixel[2:0] = 3'b000;
      14'b10110101000011: pixel[2:0] = 3'b000;
      14'b10110101000100: pixel[2:0] = 3'b000;
      14'b10110101000101: pixel[2:0] = 3'b000;
      14'b10110101000110: pixel[2:0] = 3'b000;
      14'b10110101000111: pixel[2:0] = 3'b000;
      14'b10110101001000: pixel[2:0] = 3'b000;
      14'b10110101001001: pixel[2:0] = 3'b000;
      14'b10110101001010: pixel[2:0] = 3'b000;
      14'b10110101001011: pixel[2:0] = 3'b000;
      14'b10110101001100: pixel[2:0] = 3'b000;
      14'b10110101001101: pixel[2:0] = 3'b000;
      14'b10110101001110: pixel[2:0] = 3'b000;
      14'b10110101001111: pixel[2:0] = 3'b000;
      14'b10110101010000: pixel[2:0] = 3'b000;
      14'b10110101010001: pixel[2:0] = 3'b000;
      14'b10110101010010: pixel[2:0] = 3'b000;
      14'b10110101010011: pixel[2:0] = 3'b000;
      14'b10110101010100: pixel[2:0] = 3'b000;
      14'b10110101010101: pixel[2:0] = 3'b000;
      14'b10110101010110: pixel[2:0] = 3'b000;
      14'b10110101010111: pixel[2:0] = 3'b000;
      14'b10110101011000: pixel[2:0] = 3'b000;
      14'b10110101011001: pixel[2:0] = 3'b000;
      14'b10110101011010: pixel[2:0] = 3'b000;
      14'b10110101011011: pixel[2:0] = 3'b000;
      14'b10110101011100: pixel[2:0] = 3'b000;
      14'b10110101011101: pixel[2:0] = 3'b000;
      14'b10110101011110: pixel[2:0] = 3'b000;
      14'b10110101011111: pixel[2:0] = 3'b000;
      14'b10110101100000: pixel[2:0] = 3'b000;
      14'b10110101100001: pixel[2:0] = 3'b000;
      14'b10110101100010: pixel[2:0] = 3'b000;
      14'b10110101100011: pixel[2:0] = 3'b000;
      14'b10110101100100: pixel[2:0] = 3'b000;
      14'b10110101100101: pixel[2:0] = 3'b000;
      14'b10110101100110: pixel[2:0] = 3'b000;
      14'b10110101100111: pixel[2:0] = 3'b000;
      14'b10110101101000: pixel[2:0] = 3'b000;
      14'b10110101101001: pixel[2:0] = 3'b000;
      14'b10110101101010: pixel[2:0] = 3'b000;
      14'b10110101101011: pixel[2:0] = 3'b000;
      14'b10110101101100: pixel[2:0] = 3'b000;
      14'b10110101101101: pixel[2:0] = 3'b000;
      14'b10110101101110: pixel[2:0] = 3'b000;
      14'b10110101101111: pixel[2:0] = 3'b000;
      14'b10110101110000: pixel[2:0] = 3'b000;
      14'b10110101110001: pixel[2:0] = 3'b000;
      14'b10110101110010: pixel[2:0] = 3'b000;
      14'b10110101110011: pixel[2:0] = 3'b000;
      14'b10110101110100: pixel[2:0] = 3'b000;
      14'b10110101110101: pixel[2:0] = 3'b000;
      14'b10110101110110: pixel[2:0] = 3'b000;
      14'b10110101110111: pixel[2:0] = 3'b000;
      14'b10110101111000: pixel[2:0] = 3'b000;
      14'b10110101111001: pixel[2:0] = 3'b000;
      14'b10110101111010: pixel[2:0] = 3'b000;
      14'b10110101111011: pixel[2:0] = 3'b000;
      14'b10110101111100: pixel[2:0] = 3'b000;
      14'b10110101111101: pixel[2:0] = 3'b000;
      14'b10110101111110: pixel[2:0] = 3'b000;
      14'b10110101111111: pixel[2:0] = 3'b000;
      14'b10110110000000: pixel[2:0] = 3'b000;
      14'b10110110000001: pixel[2:0] = 3'b000;
      14'b10110110000010: pixel[2:0] = 3'b000;
      14'b10110110000011: pixel[2:0] = 3'b000;
      14'b10110110000100: pixel[2:0] = 3'b000;
      14'b10110110000101: pixel[2:0] = 3'b000;
      14'b10110110000110: pixel[2:0] = 3'b000;
      14'b10110110000111: pixel[2:0] = 3'b000;
      14'b10111000000000: pixel[2:0] = 3'b000;
      14'b10111000000001: pixel[2:0] = 3'b000;
      14'b10111000000010: pixel[2:0] = 3'b000;
      14'b10111000000011: pixel[2:0] = 3'b000;
      14'b10111000000100: pixel[2:0] = 3'b000;
      14'b10111000000101: pixel[2:0] = 3'b000;
      14'b10111000000110: pixel[2:0] = 3'b000;
      14'b10111000000111: pixel[2:0] = 3'b000;
      14'b10111000001000: pixel[2:0] = 3'b000;
      14'b10111000001001: pixel[2:0] = 3'b000;
      14'b10111000001010: pixel[2:0] = 3'b000;
      14'b10111000001011: pixel[2:0] = 3'b000;
      14'b10111000001100: pixel[2:0] = 3'b000;
      14'b10111000001101: pixel[2:0] = 3'b000;
      14'b10111000001110: pixel[2:0] = 3'b000;
      14'b10111000001111: pixel[2:0] = 3'b000;
      14'b10111000010000: pixel[2:0] = 3'b000;
      14'b10111000010001: pixel[2:0] = 3'b000;
      14'b10111000010010: pixel[2:0] = 3'b000;
      14'b10111000010011: pixel[2:0] = 3'b000;
      14'b10111000010100: pixel[2:0] = 3'b000;
      14'b10111000010101: pixel[2:0] = 3'b000;
      14'b10111000010110: pixel[2:0] = 3'b000;
      14'b10111000010111: pixel[2:0] = 3'b000;
      14'b10111000011000: pixel[2:0] = 3'b000;
      14'b10111000011001: pixel[2:0] = 3'b000;
      14'b10111000011010: pixel[2:0] = 3'b000;
      14'b10111000011011: pixel[2:0] = 3'b000;
      14'b10111000011100: pixel[2:0] = 3'b000;
      14'b10111000011101: pixel[2:0] = 3'b000;
      14'b10111000011110: pixel[2:0] = 3'b000;
      14'b10111000011111: pixel[2:0] = 3'b000;
      14'b10111000100000: pixel[2:0] = 3'b000;
      14'b10111000100001: pixel[2:0] = 3'b000;
      14'b10111000100010: pixel[2:0] = 3'b000;
      14'b10111000100011: pixel[2:0] = 3'b000;
      14'b10111000100100: pixel[2:0] = 3'b000;
      14'b10111000100101: pixel[2:0] = 3'b000;
      14'b10111000100110: pixel[2:0] = 3'b000;
      14'b10111000100111: pixel[2:0] = 3'b000;
      14'b10111000101000: pixel[2:0] = 3'b000;
      14'b10111000101001: pixel[2:0] = 3'b000;
      14'b10111000101010: pixel[2:0] = 3'b000;
      14'b10111000101011: pixel[2:0] = 3'b000;
      14'b10111000101100: pixel[2:0] = 3'b000;
      14'b10111000101101: pixel[2:0] = 3'b000;
      14'b10111000101110: pixel[2:0] = 3'b000;
      14'b10111000101111: pixel[2:0] = 3'b000;
      14'b10111000110000: pixel[2:0] = 3'b000;
      14'b10111000110001: pixel[2:0] = 3'b000;
      14'b10111000110010: pixel[2:0] = 3'b000;
      14'b10111000110011: pixel[2:0] = 3'b000;
      14'b10111000110100: pixel[2:0] = 3'b000;
      14'b10111000110101: pixel[2:0] = 3'b000;
      14'b10111000110110: pixel[2:0] = 3'b000;
      14'b10111000110111: pixel[2:0] = 3'b000;
      14'b10111000111000: pixel[2:0] = 3'b000;
      14'b10111000111001: pixel[2:0] = 3'b000;
      14'b10111000111010: pixel[2:0] = 3'b000;
      14'b10111000111011: pixel[2:0] = 3'b000;
      14'b10111000111100: pixel[2:0] = 3'b000;
      14'b10111000111101: pixel[2:0] = 3'b000;
      14'b10111000111110: pixel[2:0] = 3'b000;
      14'b10111000111111: pixel[2:0] = 3'b000;
      14'b10111001000000: pixel[2:0] = 3'b000;
      14'b10111001000001: pixel[2:0] = 3'b000;
      14'b10111001000010: pixel[2:0] = 3'b000;
      14'b10111001000011: pixel[2:0] = 3'b000;
      14'b10111001000100: pixel[2:0] = 3'b000;
      14'b10111001000101: pixel[2:0] = 3'b000;
      14'b10111001000110: pixel[2:0] = 3'b000;
      14'b10111001000111: pixel[2:0] = 3'b000;
      14'b10111001001000: pixel[2:0] = 3'b000;
      14'b10111001001001: pixel[2:0] = 3'b000;
      14'b10111001001010: pixel[2:0] = 3'b000;
      14'b10111001001011: pixel[2:0] = 3'b000;
      14'b10111001001100: pixel[2:0] = 3'b000;
      14'b10111001001101: pixel[2:0] = 3'b000;
      14'b10111001001110: pixel[2:0] = 3'b000;
      14'b10111001001111: pixel[2:0] = 3'b000;
      14'b10111001010000: pixel[2:0] = 3'b000;
      14'b10111001010001: pixel[2:0] = 3'b000;
      14'b10111001010010: pixel[2:0] = 3'b000;
      14'b10111001010011: pixel[2:0] = 3'b000;
      14'b10111001010100: pixel[2:0] = 3'b000;
      14'b10111001010101: pixel[2:0] = 3'b000;
      14'b10111001010110: pixel[2:0] = 3'b000;
      14'b10111001010111: pixel[2:0] = 3'b000;
      14'b10111001011000: pixel[2:0] = 3'b000;
      14'b10111001011001: pixel[2:0] = 3'b000;
      14'b10111001011010: pixel[2:0] = 3'b000;
      14'b10111001011011: pixel[2:0] = 3'b000;
      14'b10111001011100: pixel[2:0] = 3'b000;
      14'b10111001011101: pixel[2:0] = 3'b000;
      14'b10111001011110: pixel[2:0] = 3'b000;
      14'b10111001011111: pixel[2:0] = 3'b000;
      14'b10111001100000: pixel[2:0] = 3'b000;
      14'b10111001100001: pixel[2:0] = 3'b000;
      14'b10111001100010: pixel[2:0] = 3'b000;
      14'b10111001100011: pixel[2:0] = 3'b000;
      14'b10111001100100: pixel[2:0] = 3'b000;
      14'b10111001100101: pixel[2:0] = 3'b000;
      14'b10111001100110: pixel[2:0] = 3'b000;
      14'b10111001100111: pixel[2:0] = 3'b000;
      14'b10111001101000: pixel[2:0] = 3'b000;
      14'b10111001101001: pixel[2:0] = 3'b000;
      14'b10111001101010: pixel[2:0] = 3'b000;
      14'b10111001101011: pixel[2:0] = 3'b000;
      14'b10111001101100: pixel[2:0] = 3'b000;
      14'b10111001101101: pixel[2:0] = 3'b000;
      14'b10111001101110: pixel[2:0] = 3'b000;
      14'b10111001101111: pixel[2:0] = 3'b000;
      14'b10111001110000: pixel[2:0] = 3'b000;
      14'b10111001110001: pixel[2:0] = 3'b000;
      14'b10111001110010: pixel[2:0] = 3'b000;
      14'b10111001110011: pixel[2:0] = 3'b000;
      14'b10111001110100: pixel[2:0] = 3'b000;
      14'b10111001110101: pixel[2:0] = 3'b000;
      14'b10111001110110: pixel[2:0] = 3'b000;
      14'b10111001110111: pixel[2:0] = 3'b000;
      14'b10111001111000: pixel[2:0] = 3'b000;
      14'b10111001111001: pixel[2:0] = 3'b000;
      14'b10111001111010: pixel[2:0] = 3'b000;
      14'b10111001111011: pixel[2:0] = 3'b000;
      14'b10111001111100: pixel[2:0] = 3'b000;
      14'b10111001111101: pixel[2:0] = 3'b000;
      14'b10111001111110: pixel[2:0] = 3'b000;
      14'b10111001111111: pixel[2:0] = 3'b000;
      14'b10111010000000: pixel[2:0] = 3'b000;
      14'b10111010000001: pixel[2:0] = 3'b000;
      14'b10111010000010: pixel[2:0] = 3'b000;
      14'b10111010000011: pixel[2:0] = 3'b000;
      14'b10111010000100: pixel[2:0] = 3'b000;
      14'b10111010000101: pixel[2:0] = 3'b000;
      14'b10111010000110: pixel[2:0] = 3'b000;
      14'b10111010000111: pixel[2:0] = 3'b000;
      14'b10111100000000: pixel[2:0] = 3'b000;
      14'b10111100000001: pixel[2:0] = 3'b000;
      14'b10111100000010: pixel[2:0] = 3'b000;
      14'b10111100000011: pixel[2:0] = 3'b000;
      14'b10111100000100: pixel[2:0] = 3'b000;
      14'b10111100000101: pixel[2:0] = 3'b000;
      14'b10111100000110: pixel[2:0] = 3'b000;
      14'b10111100000111: pixel[2:0] = 3'b000;
      14'b10111100001000: pixel[2:0] = 3'b000;
      14'b10111100001001: pixel[2:0] = 3'b000;
      14'b10111100001010: pixel[2:0] = 3'b000;
      14'b10111100001011: pixel[2:0] = 3'b000;
      14'b10111100001100: pixel[2:0] = 3'b000;
      14'b10111100001101: pixel[2:0] = 3'b000;
      14'b10111100001110: pixel[2:0] = 3'b000;
      14'b10111100001111: pixel[2:0] = 3'b000;
      14'b10111100010000: pixel[2:0] = 3'b000;
      14'b10111100010001: pixel[2:0] = 3'b000;
      14'b10111100010010: pixel[2:0] = 3'b000;
      14'b10111100010011: pixel[2:0] = 3'b000;
      14'b10111100010100: pixel[2:0] = 3'b000;
      14'b10111100010101: pixel[2:0] = 3'b000;
      14'b10111100010110: pixel[2:0] = 3'b000;
      14'b10111100010111: pixel[2:0] = 3'b000;
      14'b10111100011000: pixel[2:0] = 3'b000;
      14'b10111100011001: pixel[2:0] = 3'b000;
      14'b10111100011010: pixel[2:0] = 3'b000;
      14'b10111100011011: pixel[2:0] = 3'b000;
      14'b10111100011100: pixel[2:0] = 3'b000;
      14'b10111100011101: pixel[2:0] = 3'b000;
      14'b10111100011110: pixel[2:0] = 3'b000;
      14'b10111100011111: pixel[2:0] = 3'b000;
      14'b10111100100000: pixel[2:0] = 3'b000;
      14'b10111100100001: pixel[2:0] = 3'b000;
      14'b10111100100010: pixel[2:0] = 3'b000;
      14'b10111100100011: pixel[2:0] = 3'b000;
      14'b10111100100100: pixel[2:0] = 3'b000;
      14'b10111100100101: pixel[2:0] = 3'b000;
      14'b10111100100110: pixel[2:0] = 3'b000;
      14'b10111100100111: pixel[2:0] = 3'b000;
      14'b10111100101000: pixel[2:0] = 3'b000;
      14'b10111100101001: pixel[2:0] = 3'b000;
      14'b10111100101010: pixel[2:0] = 3'b000;
      14'b10111100101011: pixel[2:0] = 3'b000;
      14'b10111100101100: pixel[2:0] = 3'b000;
      14'b10111100101101: pixel[2:0] = 3'b000;
      14'b10111100101110: pixel[2:0] = 3'b000;
      14'b10111100101111: pixel[2:0] = 3'b000;
      14'b10111100110000: pixel[2:0] = 3'b000;
      14'b10111100110001: pixel[2:0] = 3'b000;
      14'b10111100110010: pixel[2:0] = 3'b000;
      14'b10111100110011: pixel[2:0] = 3'b000;
      14'b10111100110100: pixel[2:0] = 3'b000;
      14'b10111100110101: pixel[2:0] = 3'b000;
      14'b10111100110110: pixel[2:0] = 3'b000;
      14'b10111100110111: pixel[2:0] = 3'b000;
      14'b10111100111000: pixel[2:0] = 3'b000;
      14'b10111100111001: pixel[2:0] = 3'b000;
      14'b10111100111010: pixel[2:0] = 3'b000;
      14'b10111100111011: pixel[2:0] = 3'b000;
      14'b10111100111100: pixel[2:0] = 3'b000;
      14'b10111100111101: pixel[2:0] = 3'b000;
      14'b10111100111110: pixel[2:0] = 3'b000;
      14'b10111100111111: pixel[2:0] = 3'b000;
      14'b10111101000000: pixel[2:0] = 3'b000;
      14'b10111101000001: pixel[2:0] = 3'b000;
      14'b10111101000010: pixel[2:0] = 3'b000;
      14'b10111101000011: pixel[2:0] = 3'b000;
      14'b10111101000100: pixel[2:0] = 3'b000;
      14'b10111101000101: pixel[2:0] = 3'b000;
      14'b10111101000110: pixel[2:0] = 3'b000;
      14'b10111101000111: pixel[2:0] = 3'b000;
      14'b10111101001000: pixel[2:0] = 3'b000;
      14'b10111101001001: pixel[2:0] = 3'b000;
      14'b10111101001010: pixel[2:0] = 3'b000;
      14'b10111101001011: pixel[2:0] = 3'b000;
      14'b10111101001100: pixel[2:0] = 3'b000;
      14'b10111101001101: pixel[2:0] = 3'b000;
      14'b10111101001110: pixel[2:0] = 3'b000;
      14'b10111101001111: pixel[2:0] = 3'b000;
      14'b10111101010000: pixel[2:0] = 3'b000;
      14'b10111101010001: pixel[2:0] = 3'b000;
      14'b10111101010010: pixel[2:0] = 3'b000;
      14'b10111101010011: pixel[2:0] = 3'b000;
      14'b10111101010100: pixel[2:0] = 3'b000;
      14'b10111101010101: pixel[2:0] = 3'b000;
      14'b10111101010110: pixel[2:0] = 3'b000;
      14'b10111101010111: pixel[2:0] = 3'b000;
      14'b10111101011000: pixel[2:0] = 3'b000;
      14'b10111101011001: pixel[2:0] = 3'b000;
      14'b10111101011010: pixel[2:0] = 3'b000;
      14'b10111101011011: pixel[2:0] = 3'b000;
      14'b10111101011100: pixel[2:0] = 3'b000;
      14'b10111101011101: pixel[2:0] = 3'b000;
      14'b10111101011110: pixel[2:0] = 3'b000;
      14'b10111101011111: pixel[2:0] = 3'b000;
      14'b10111101100000: pixel[2:0] = 3'b000;
      14'b10111101100001: pixel[2:0] = 3'b000;
      14'b10111101100010: pixel[2:0] = 3'b000;
      14'b10111101100011: pixel[2:0] = 3'b000;
      14'b10111101100100: pixel[2:0] = 3'b000;
      14'b10111101100101: pixel[2:0] = 3'b000;
      14'b10111101100110: pixel[2:0] = 3'b000;
      14'b10111101100111: pixel[2:0] = 3'b000;
      14'b10111101101000: pixel[2:0] = 3'b000;
      14'b10111101101001: pixel[2:0] = 3'b000;
      14'b10111101101010: pixel[2:0] = 3'b000;
      14'b10111101101011: pixel[2:0] = 3'b000;
      14'b10111101101100: pixel[2:0] = 3'b000;
      14'b10111101101101: pixel[2:0] = 3'b000;
      14'b10111101101110: pixel[2:0] = 3'b000;
      14'b10111101101111: pixel[2:0] = 3'b000;
      14'b10111101110000: pixel[2:0] = 3'b000;
      14'b10111101110001: pixel[2:0] = 3'b000;
      14'b10111101110010: pixel[2:0] = 3'b000;
      14'b10111101110011: pixel[2:0] = 3'b000;
      14'b10111101110100: pixel[2:0] = 3'b000;
      14'b10111101110101: pixel[2:0] = 3'b000;
      14'b10111101110110: pixel[2:0] = 3'b000;
      14'b10111101110111: pixel[2:0] = 3'b000;
      14'b10111101111000: pixel[2:0] = 3'b000;
      14'b10111101111001: pixel[2:0] = 3'b000;
      14'b10111101111010: pixel[2:0] = 3'b000;
      14'b10111101111011: pixel[2:0] = 3'b000;
      14'b10111101111100: pixel[2:0] = 3'b000;
      14'b10111101111101: pixel[2:0] = 3'b000;
      14'b10111101111110: pixel[2:0] = 3'b000;
      14'b10111101111111: pixel[2:0] = 3'b000;
      14'b10111110000000: pixel[2:0] = 3'b000;
      14'b10111110000001: pixel[2:0] = 3'b000;
      14'b10111110000010: pixel[2:0] = 3'b000;
      14'b10111110000011: pixel[2:0] = 3'b000;
      14'b10111110000100: pixel[2:0] = 3'b000;
      14'b10111110000101: pixel[2:0] = 3'b000;
      14'b10111110000110: pixel[2:0] = 3'b000;
      14'b10111110000111: pixel[2:0] = 3'b000;
    default: pixel = 3'b000;
  endcase
endmodule
